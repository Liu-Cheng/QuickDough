`timescale 1ns / 1ps

module torus100(
	      clk,
          rst_n,
          data_out0,
          data_out1,
          data_out2,
          data_out3
	      );

input clk;
input rst_n;

output[15:0] data_out0;
output[15:0] data_out1;
output[15:0] data_out2;
output[15:0] data_out3;

wire [15:0] PE00_out0;
wire [15:0] PE00_out1;
wire [15:0] PE00_out2;
wire [15:0] PE00_out3;

wire [15:0] PE01_out0;
wire [15:0] PE01_out1;
wire [15:0] PE01_out2;
wire [15:0] PE01_out3;

wire [15:0] PE02_out0;
wire [15:0] PE02_out1;
wire [15:0] PE02_out2;
wire [15:0] PE02_out3;

wire [15:0] PE03_out0;
wire [15:0] PE03_out1;
wire [15:0] PE03_out2;
wire [15:0] PE03_out3;

wire [15:0] PE04_out0;
wire [15:0] PE04_out1;
wire [15:0] PE04_out2;
wire [15:0] PE04_out3;

wire [15:0] PE05_out0;
wire [15:0] PE05_out1;
wire [15:0] PE05_out2;
wire [15:0] PE05_out3;

wire [15:0] PE06_out0;
wire [15:0] PE06_out1;
wire [15:0] PE06_out2;
wire [15:0] PE06_out3;

wire [15:0] PE07_out0;
wire [15:0] PE07_out1;
wire [15:0] PE07_out2;
wire [15:0] PE07_out3;

wire [15:0] PE08_out0;
wire [15:0] PE08_out1;
wire [15:0] PE08_out2;
wire [15:0] PE08_out3;

wire [15:0] PE09_out0;
wire [15:0] PE09_out1;
wire [15:0] PE09_out2;
wire [15:0] PE09_out3;


wire [15:0] PE10_out0;
wire [15:0] PE10_out1;
wire [15:0] PE10_out2;
wire [15:0] PE10_out3;

wire [15:0] PE11_out0;
wire [15:0] PE11_out1;
wire [15:0] PE11_out2;
wire [15:0] PE11_out3;

wire [15:0] PE12_out0;
wire [15:0] PE12_out1;
wire [15:0] PE12_out2;
wire [15:0] PE12_out3;

wire [15:0] PE13_out0;
wire [15:0] PE13_out1;
wire [15:0] PE13_out2;
wire [15:0] PE13_out3;

wire [15:0] PE14_out0;
wire [15:0] PE14_out1;
wire [15:0] PE14_out2;
wire [15:0] PE14_out3;

wire [15:0] PE15_out0;
wire [15:0] PE15_out1;
wire [15:0] PE15_out2;
wire [15:0] PE15_out3;

wire [15:0] PE16_out0;
wire [15:0] PE16_out1;
wire [15:0] PE16_out2;
wire [15:0] PE16_out3;

wire [15:0] PE17_out0;
wire [15:0] PE17_out1;
wire [15:0] PE17_out2;
wire [15:0] PE17_out3;

wire [15:0] PE18_out0;
wire [15:0] PE18_out1;
wire [15:0] PE18_out2;
wire [15:0] PE18_out3;

wire [15:0] PE19_out0;
wire [15:0] PE19_out1;
wire [15:0] PE19_out2;
wire [15:0] PE19_out3;


wire [15:0] PE20_out0;
wire [15:0] PE20_out1;
wire [15:0] PE20_out2;
wire [15:0] PE20_out3;

wire [15:0] PE21_out0;
wire [15:0] PE21_out1;
wire [15:0] PE21_out2;
wire [15:0] PE21_out3;

wire [15:0] PE22_out0;
wire [15:0] PE22_out1;
wire [15:0] PE22_out2;
wire [15:0] PE22_out3;

wire [15:0] PE23_out0;
wire [15:0] PE23_out1;
wire [15:0] PE23_out2;
wire [15:0] PE23_out3;

wire [15:0] PE24_out0;
wire [15:0] PE24_out1;
wire [15:0] PE24_out2;
wire [15:0] PE24_out3;

wire [15:0] PE25_out0;
wire [15:0] PE25_out1;
wire [15:0] PE25_out2;
wire [15:0] PE25_out3;

wire [15:0] PE26_out0;
wire [15:0] PE26_out1;
wire [15:0] PE26_out2;
wire [15:0] PE26_out3;

wire [15:0] PE27_out0;
wire [15:0] PE27_out1;
wire [15:0] PE27_out2;
wire [15:0] PE27_out3;

wire [15:0] PE28_out0;
wire [15:0] PE28_out1;
wire [15:0] PE28_out2;
wire [15:0] PE28_out3;

wire [15:0] PE29_out0;
wire [15:0] PE29_out1;
wire [15:0] PE29_out2;
wire [15:0] PE29_out3;


wire [15:0] PE30_out0;
wire [15:0] PE30_out1;
wire [15:0] PE30_out2;
wire [15:0] PE30_out3;

wire [15:0] PE31_out0;
wire [15:0] PE31_out1;
wire [15:0] PE31_out2;
wire [15:0] PE31_out3;

wire [15:0] PE32_out0;
wire [15:0] PE32_out1;
wire [15:0] PE32_out2;
wire [15:0] PE32_out3;

wire [15:0] PE33_out0;
wire [15:0] PE33_out1;
wire [15:0] PE33_out2;
wire [15:0] PE33_out3;

wire [15:0] PE34_out0;
wire [15:0] PE34_out1;
wire [15:0] PE34_out2;
wire [15:0] PE34_out3;

wire [15:0] PE35_out0;
wire [15:0] PE35_out1;
wire [15:0] PE35_out2;
wire [15:0] PE35_out3;

wire [15:0] PE36_out0;
wire [15:0] PE36_out1;
wire [15:0] PE36_out2;
wire [15:0] PE36_out3;

wire [15:0] PE37_out0;
wire [15:0] PE37_out1;
wire [15:0] PE37_out2;
wire [15:0] PE37_out3;

wire [15:0] PE38_out0;
wire [15:0] PE38_out1;
wire [15:0] PE38_out2;
wire [15:0] PE38_out3;

wire [15:0] PE39_out0;
wire [15:0] PE39_out1;
wire [15:0] PE39_out2;
wire [15:0] PE39_out3;


wire [15:0] PE40_out0;
wire [15:0] PE40_out1;
wire [15:0] PE40_out2;
wire [15:0] PE40_out3;

wire [15:0] PE41_out0;
wire [15:0] PE41_out1;
wire [15:0] PE41_out2;
wire [15:0] PE41_out3;

wire [15:0] PE42_out0;
wire [15:0] PE42_out1;
wire [15:0] PE42_out2;
wire [15:0] PE42_out3;

wire [15:0] PE43_out0;
wire [15:0] PE43_out1;
wire [15:0] PE43_out2;
wire [15:0] PE43_out3;

wire [15:0] PE44_out0;
wire [15:0] PE44_out1;
wire [15:0] PE44_out2;
wire [15:0] PE44_out3;

wire [15:0] PE45_out0;
wire [15:0] PE45_out1;
wire [15:0] PE45_out2;
wire [15:0] PE45_out3;

wire [15:0] PE46_out0;
wire [15:0] PE46_out1;
wire [15:0] PE46_out2;
wire [15:0] PE46_out3;

wire [15:0] PE47_out0;
wire [15:0] PE47_out1;
wire [15:0] PE47_out2;
wire [15:0] PE47_out3;

wire [15:0] PE48_out0;
wire [15:0] PE48_out1;
wire [15:0] PE48_out2;
wire [15:0] PE48_out3;

wire [15:0] PE49_out0;
wire [15:0] PE49_out1;
wire [15:0] PE49_out2;
wire [15:0] PE49_out3;


wire [15:0] PE50_out0;
wire [15:0] PE50_out1;
wire [15:0] PE50_out2;
wire [15:0] PE50_out3;

wire [15:0] PE51_out0;
wire [15:0] PE51_out1;
wire [15:0] PE51_out2;
wire [15:0] PE51_out3;

wire [15:0] PE52_out0;
wire [15:0] PE52_out1;
wire [15:0] PE52_out2;
wire [15:0] PE52_out3;

wire [15:0] PE53_out0;
wire [15:0] PE53_out1;
wire [15:0] PE53_out2;
wire [15:0] PE53_out3;

wire [15:0] PE54_out0;
wire [15:0] PE54_out1;
wire [15:0] PE54_out2;
wire [15:0] PE54_out3;

wire [15:0] PE55_out0;
wire [15:0] PE55_out1;
wire [15:0] PE55_out2;
wire [15:0] PE55_out3;

wire [15:0] PE56_out0;
wire [15:0] PE56_out1;
wire [15:0] PE56_out2;
wire [15:0] PE56_out3;

wire [15:0] PE57_out0;
wire [15:0] PE57_out1;
wire [15:0] PE57_out2;
wire [15:0] PE57_out3;

wire [15:0] PE58_out0;
wire [15:0] PE58_out1;
wire [15:0] PE58_out2;
wire [15:0] PE58_out3;

wire [15:0] PE59_out0;
wire [15:0] PE59_out1;
wire [15:0] PE59_out2;
wire [15:0] PE59_out3;


wire [15:0] PE60_out0;
wire [15:0] PE60_out1;
wire [15:0] PE60_out2;
wire [15:0] PE60_out3;

wire [15:0] PE61_out0;
wire [15:0] PE61_out1;
wire [15:0] PE61_out2;
wire [15:0] PE61_out3;

wire [15:0] PE62_out0;
wire [15:0] PE62_out1;
wire [15:0] PE62_out2;
wire [15:0] PE62_out3;

wire [15:0] PE63_out0;
wire [15:0] PE63_out1;
wire [15:0] PE63_out2;
wire [15:0] PE63_out3;

wire [15:0] PE64_out0;
wire [15:0] PE64_out1;
wire [15:0] PE64_out2;
wire [15:0] PE64_out3;

wire [15:0] PE65_out0;
wire [15:0] PE65_out1;
wire [15:0] PE65_out2;
wire [15:0] PE65_out3;

wire [15:0] PE66_out0;
wire [15:0] PE66_out1;
wire [15:0] PE66_out2;
wire [15:0] PE66_out3;

wire [15:0] PE67_out0;
wire [15:0] PE67_out1;
wire [15:0] PE67_out2;
wire [15:0] PE67_out3;

wire [15:0] PE68_out0;
wire [15:0] PE68_out1;
wire [15:0] PE68_out2;
wire [15:0] PE68_out3;

wire [15:0] PE69_out0;
wire [15:0] PE69_out1;
wire [15:0] PE69_out2;
wire [15:0] PE69_out3;


wire [15:0] PE70_out0;
wire [15:0] PE70_out1;
wire [15:0] PE70_out2;
wire [15:0] PE70_out3;

wire [15:0] PE71_out0;
wire [15:0] PE71_out1;
wire [15:0] PE71_out2;
wire [15:0] PE71_out3;

wire [15:0] PE72_out0;
wire [15:0] PE72_out1;
wire [15:0] PE72_out2;
wire [15:0] PE72_out3;

wire [15:0] PE73_out0;
wire [15:0] PE73_out1;
wire [15:0] PE73_out2;
wire [15:0] PE73_out3;

wire [15:0] PE74_out0;
wire [15:0] PE74_out1;
wire [15:0] PE74_out2;
wire [15:0] PE74_out3;

wire [15:0] PE75_out0;
wire [15:0] PE75_out1;
wire [15:0] PE75_out2;
wire [15:0] PE75_out3;

wire [15:0] PE76_out0;
wire [15:0] PE76_out1;
wire [15:0] PE76_out2;
wire [15:0] PE76_out3;

wire [15:0] PE77_out0;
wire [15:0] PE77_out1;
wire [15:0] PE77_out2;
wire [15:0] PE77_out3;

wire [15:0] PE78_out0;
wire [15:0] PE78_out1;
wire [15:0] PE78_out2;
wire [15:0] PE78_out3;

wire [15:0] PE79_out0;
wire [15:0] PE79_out1;
wire [15:0] PE79_out2;
wire [15:0] PE79_out3;


wire [15:0] PE80_out0;
wire [15:0] PE80_out1;
wire [15:0] PE80_out2;
wire [15:0] PE80_out3;

wire [15:0] PE81_out0;
wire [15:0] PE81_out1;
wire [15:0] PE81_out2;
wire [15:0] PE81_out3;

wire [15:0] PE82_out0;
wire [15:0] PE82_out1;
wire [15:0] PE82_out2;
wire [15:0] PE82_out3;

wire [15:0] PE83_out0;
wire [15:0] PE83_out1;
wire [15:0] PE83_out2;
wire [15:0] PE83_out3;

wire [15:0] PE84_out0;
wire [15:0] PE84_out1;
wire [15:0] PE84_out2;
wire [15:0] PE84_out3;

wire [15:0] PE85_out0;
wire [15:0] PE85_out1;
wire [15:0] PE85_out2;
wire [15:0] PE85_out3;

wire [15:0] PE86_out0;
wire [15:0] PE86_out1;
wire [15:0] PE86_out2;
wire [15:0] PE86_out3;

wire [15:0] PE87_out0;
wire [15:0] PE87_out1;
wire [15:0] PE87_out2;
wire [15:0] PE87_out3;

wire [15:0] PE88_out0;
wire [15:0] PE88_out1;
wire [15:0] PE88_out2;
wire [15:0] PE88_out3;

wire [15:0] PE89_out0;
wire [15:0] PE89_out1;
wire [15:0] PE89_out2;
wire [15:0] PE89_out3;


wire [15:0] PE90_out0;
wire [15:0] PE90_out1;
wire [15:0] PE90_out2;
wire [15:0] PE90_out3;

wire [15:0] PE91_out0;
wire [15:0] PE91_out1;
wire [15:0] PE91_out2;
wire [15:0] PE91_out3;

wire [15:0] PE92_out0;
wire [15:0] PE92_out1;
wire [15:0] PE92_out2;
wire [15:0] PE92_out3;

wire [15:0] PE93_out0;
wire [15:0] PE93_out1;
wire [15:0] PE93_out2;
wire [15:0] PE93_out3;

wire [15:0] PE94_out0;
wire [15:0] PE94_out1;
wire [15:0] PE94_out2;
wire [15:0] PE94_out3;

wire [15:0] PE95_out0;
wire [15:0] PE95_out1;
wire [15:0] PE95_out2;
wire [15:0] PE95_out3;

wire [15:0] PE96_out0;
wire [15:0] PE96_out1;
wire [15:0] PE96_out2;
wire [15:0] PE96_out3;

wire [15:0] PE97_out0;
wire [15:0] PE97_out1;
wire [15:0] PE97_out2;
wire [15:0] PE97_out3;

wire [15:0] PE98_out0;
wire [15:0] PE98_out1;
wire [15:0] PE98_out2;
wire [15:0] PE98_out3;

wire [15:0] PE99_out0;
wire [15:0] PE99_out1;
wire [15:0] PE99_out2;
wire [15:0] PE99_out3;



PE PE00(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE09_out2),
     .PE_in1(PE90_out3),
     .PE_in2(PE01_out0),
     .PE_in3(PE10_out1),

     .PE_out0(PE00_out0),
     .PE_out1(PE00_out1),
     .PE_out2(PE00_out2),
     .PE_out3(PE00_out3)
       );

PE PE01(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE00_out2),
     .PE_in1(PE91_out3),
     .PE_in2(PE02_out0),
     .PE_in3(PE11_out1),

     .PE_out0(PE01_out0),
     .PE_out1(PE01_out1),
     .PE_out2(PE01_out2),
     .PE_out3(PE01_out3)
       );

PE PE02(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE01_out2),
     .PE_in1(PE92_out3),
     .PE_in2(PE03_out0),
     .PE_in3(PE12_out1),

     .PE_out0(PE02_out0),
     .PE_out1(PE02_out1),
     .PE_out2(PE02_out2),
     .PE_out3(PE02_out3)
       );

PE PE03(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE02_out2),
     .PE_in1(PE93_out3),
     .PE_in2(PE04_out0),
     .PE_in3(PE13_out1),

     .PE_out0(PE03_out0),
     .PE_out1(PE03_out1),
     .PE_out2(PE03_out2),
     .PE_out3(PE03_out3)
       );

PE PE04(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE03_out2),
     .PE_in1(PE94_out3),
     .PE_in2(PE05_out0),
     .PE_in3(PE14_out1),

     .PE_out0(PE04_out0),
     .PE_out1(PE04_out1),
     .PE_out2(PE04_out2),
     .PE_out3(PE04_out3)
       );

PE PE05(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE04_out2),
     .PE_in1(PE95_out3),
     .PE_in2(PE06_out0),
     .PE_in3(PE15_out1),

     .PE_out0(PE05_out0),
     .PE_out1(PE05_out1),
     .PE_out2(PE05_out2),
     .PE_out3(PE05_out3)
       );

PE PE06(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE05_out2),
     .PE_in1(PE96_out3),
     .PE_in2(PE07_out0),
     .PE_in3(PE16_out1),

     .PE_out0(PE06_out0),
     .PE_out1(PE06_out1),
     .PE_out2(PE06_out2),
     .PE_out3(PE06_out3)
       );

PE PE07(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE06_out2),
     .PE_in1(PE97_out3),
     .PE_in2(PE08_out0),
     .PE_in3(PE17_out1),

     .PE_out0(PE07_out0),
     .PE_out1(PE07_out1),
     .PE_out2(PE07_out2),
     .PE_out3(PE07_out3)
       );

PE PE08(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE07_out2),
     .PE_in1(PE98_out3),
     .PE_in2(PE09_out0),
     .PE_in3(PE18_out1),

     .PE_out0(PE08_out0),
     .PE_out1(PE08_out1),
     .PE_out2(PE08_out2),
     .PE_out3(PE08_out3)
       );

PE PE09(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE08_out2),
     .PE_in1(PE99_out3),
     .PE_in2(PE00_out0),
     .PE_in3(PE19_out1),

     .PE_out0(PE09_out0),
     .PE_out1(PE09_out1),
     .PE_out2(PE09_out2),
     .PE_out3(PE09_out3)
       );


PE PE10(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE19_out2),
     .PE_in1(PE00_out3),
     .PE_in2(PE11_out0),
     .PE_in3(PE20_out1),

     .PE_out0(PE10_out0),
     .PE_out1(PE10_out1),
     .PE_out2(PE10_out2),
     .PE_out3(PE10_out3)
       );

PE PE11(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE10_out2),
     .PE_in1(PE01_out3),
     .PE_in2(PE12_out0),
     .PE_in3(PE21_out1),

     .PE_out0(PE11_out0),
     .PE_out1(PE11_out1),
     .PE_out2(PE11_out2),
     .PE_out3(PE11_out3)
       );

PE PE12(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE11_out2),
     .PE_in1(PE02_out3),
     .PE_in2(PE13_out0),
     .PE_in3(PE22_out1),

     .PE_out0(PE12_out0),
     .PE_out1(PE12_out1),
     .PE_out2(PE12_out2),
     .PE_out3(PE12_out3)
       );

PE PE13(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE12_out2),
     .PE_in1(PE03_out3),
     .PE_in2(PE14_out0),
     .PE_in3(PE23_out1),

     .PE_out0(PE13_out0),
     .PE_out1(PE13_out1),
     .PE_out2(PE13_out2),
     .PE_out3(PE13_out3)
       );

PE PE14(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE13_out2),
     .PE_in1(PE04_out3),
     .PE_in2(PE15_out0),
     .PE_in3(PE24_out1),

     .PE_out0(PE14_out0),
     .PE_out1(PE14_out1),
     .PE_out2(PE14_out2),
     .PE_out3(PE14_out3)
       );

PE PE15(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE14_out2),
     .PE_in1(PE05_out3),
     .PE_in2(PE16_out0),
     .PE_in3(PE25_out1),

     .PE_out0(PE15_out0),
     .PE_out1(PE15_out1),
     .PE_out2(PE15_out2),
     .PE_out3(PE15_out3)
       );

PE PE16(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE15_out2),
     .PE_in1(PE06_out3),
     .PE_in2(PE17_out0),
     .PE_in3(PE26_out1),

     .PE_out0(PE16_out0),
     .PE_out1(PE16_out1),
     .PE_out2(PE16_out2),
     .PE_out3(PE16_out3)
       );

PE PE17(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE16_out2),
     .PE_in1(PE07_out3),
     .PE_in2(PE18_out0),
     .PE_in3(PE27_out1),

     .PE_out0(PE17_out0),
     .PE_out1(PE17_out1),
     .PE_out2(PE17_out2),
     .PE_out3(PE17_out3)
       );

PE PE18(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE17_out2),
     .PE_in1(PE08_out3),
     .PE_in2(PE19_out0),
     .PE_in3(PE28_out1),

     .PE_out0(PE18_out0),
     .PE_out1(PE18_out1),
     .PE_out2(PE18_out2),
     .PE_out3(PE18_out3)
       );

PE PE19(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE18_out2),
     .PE_in1(PE09_out3),
     .PE_in2(PE10_out0),
     .PE_in3(PE29_out1),

     .PE_out0(PE19_out0),
     .PE_out1(PE19_out1),
     .PE_out2(PE19_out2),
     .PE_out3(PE19_out3)
       );


PE PE20(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE29_out2),
     .PE_in1(PE10_out3),
     .PE_in2(PE21_out0),
     .PE_in3(PE30_out1),

     .PE_out0(PE20_out0),
     .PE_out1(PE20_out1),
     .PE_out2(PE20_out2),
     .PE_out3(PE20_out3)
       );

PE PE21(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE20_out2),
     .PE_in1(PE11_out3),
     .PE_in2(PE22_out0),
     .PE_in3(PE31_out1),

     .PE_out0(PE21_out0),
     .PE_out1(PE21_out1),
     .PE_out2(PE21_out2),
     .PE_out3(PE21_out3)
       );

PE PE22(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE21_out2),
     .PE_in1(PE12_out3),
     .PE_in2(PE23_out0),
     .PE_in3(PE32_out1),

     .PE_out0(PE22_out0),
     .PE_out1(PE22_out1),
     .PE_out2(PE22_out2),
     .PE_out3(PE22_out3)
       );

PE PE23(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE22_out2),
     .PE_in1(PE13_out3),
     .PE_in2(PE24_out0),
     .PE_in3(PE33_out1),

     .PE_out0(PE23_out0),
     .PE_out1(PE23_out1),
     .PE_out2(PE23_out2),
     .PE_out3(PE23_out3)
       );

PE PE24(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE23_out2),
     .PE_in1(PE14_out3),
     .PE_in2(PE25_out0),
     .PE_in3(PE34_out1),

     .PE_out0(PE24_out0),
     .PE_out1(PE24_out1),
     .PE_out2(PE24_out2),
     .PE_out3(PE24_out3)
       );

PE PE25(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE24_out2),
     .PE_in1(PE15_out3),
     .PE_in2(PE26_out0),
     .PE_in3(PE35_out1),

     .PE_out0(PE25_out0),
     .PE_out1(PE25_out1),
     .PE_out2(PE25_out2),
     .PE_out3(PE25_out3)
       );

PE PE26(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE25_out2),
     .PE_in1(PE16_out3),
     .PE_in2(PE27_out0),
     .PE_in3(PE36_out1),

     .PE_out0(PE26_out0),
     .PE_out1(PE26_out1),
     .PE_out2(PE26_out2),
     .PE_out3(PE26_out3)
       );

PE PE27(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE26_out2),
     .PE_in1(PE17_out3),
     .PE_in2(PE28_out0),
     .PE_in3(PE37_out1),

     .PE_out0(PE27_out0),
     .PE_out1(PE27_out1),
     .PE_out2(PE27_out2),
     .PE_out3(PE27_out3)
       );

PE PE28(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE27_out2),
     .PE_in1(PE18_out3),
     .PE_in2(PE29_out0),
     .PE_in3(PE38_out1),

     .PE_out0(PE28_out0),
     .PE_out1(PE28_out1),
     .PE_out2(PE28_out2),
     .PE_out3(PE28_out3)
       );

PE PE29(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE28_out2),
     .PE_in1(PE19_out3),
     .PE_in2(PE20_out0),
     .PE_in3(PE39_out1),

     .PE_out0(PE29_out0),
     .PE_out1(PE29_out1),
     .PE_out2(PE29_out2),
     .PE_out3(PE29_out3)
       );


PE PE30(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE39_out2),
     .PE_in1(PE20_out3),
     .PE_in2(PE31_out0),
     .PE_in3(PE40_out1),

     .PE_out0(PE30_out0),
     .PE_out1(PE30_out1),
     .PE_out2(PE30_out2),
     .PE_out3(PE30_out3)
       );

PE PE31(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE30_out2),
     .PE_in1(PE21_out3),
     .PE_in2(PE32_out0),
     .PE_in3(PE41_out1),

     .PE_out0(PE31_out0),
     .PE_out1(PE31_out1),
     .PE_out2(PE31_out2),
     .PE_out3(PE31_out3)
       );

PE PE32(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE31_out2),
     .PE_in1(PE22_out3),
     .PE_in2(PE33_out0),
     .PE_in3(PE42_out1),

     .PE_out0(PE32_out0),
     .PE_out1(PE32_out1),
     .PE_out2(PE32_out2),
     .PE_out3(PE32_out3)
       );

PE PE33(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE32_out2),
     .PE_in1(PE23_out3),
     .PE_in2(PE34_out0),
     .PE_in3(PE43_out1),

     .PE_out0(PE33_out0),
     .PE_out1(PE33_out1),
     .PE_out2(PE33_out2),
     .PE_out3(PE33_out3)
       );

PE PE34(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE33_out2),
     .PE_in1(PE24_out3),
     .PE_in2(PE35_out0),
     .PE_in3(PE44_out1),

     .PE_out0(PE34_out0),
     .PE_out1(PE34_out1),
     .PE_out2(PE34_out2),
     .PE_out3(PE34_out3)
       );

PE PE35(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE34_out2),
     .PE_in1(PE25_out3),
     .PE_in2(PE36_out0),
     .PE_in3(PE45_out1),

     .PE_out0(PE35_out0),
     .PE_out1(PE35_out1),
     .PE_out2(PE35_out2),
     .PE_out3(PE35_out3)
       );

PE PE36(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE35_out2),
     .PE_in1(PE26_out3),
     .PE_in2(PE37_out0),
     .PE_in3(PE46_out1),

     .PE_out0(PE36_out0),
     .PE_out1(PE36_out1),
     .PE_out2(PE36_out2),
     .PE_out3(PE36_out3)
       );

PE PE37(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE36_out2),
     .PE_in1(PE27_out3),
     .PE_in2(PE38_out0),
     .PE_in3(PE47_out1),

     .PE_out0(PE37_out0),
     .PE_out1(PE37_out1),
     .PE_out2(PE37_out2),
     .PE_out3(PE37_out3)
       );

PE PE38(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE37_out2),
     .PE_in1(PE28_out3),
     .PE_in2(PE39_out0),
     .PE_in3(PE48_out1),

     .PE_out0(PE38_out0),
     .PE_out1(PE38_out1),
     .PE_out2(PE38_out2),
     .PE_out3(PE38_out3)
       );

PE PE39(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE38_out2),
     .PE_in1(PE29_out3),
     .PE_in2(PE30_out0),
     .PE_in3(PE49_out1),

     .PE_out0(PE39_out0),
     .PE_out1(PE39_out1),
     .PE_out2(PE39_out2),
     .PE_out3(PE39_out3)
       );


PE PE40(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE49_out2),
     .PE_in1(PE30_out3),
     .PE_in2(PE41_out0),
     .PE_in3(PE50_out1),

     .PE_out0(PE40_out0),
     .PE_out1(PE40_out1),
     .PE_out2(PE40_out2),
     .PE_out3(PE40_out3)
       );

PE PE41(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE40_out2),
     .PE_in1(PE31_out3),
     .PE_in2(PE42_out0),
     .PE_in3(PE51_out1),

     .PE_out0(PE41_out0),
     .PE_out1(PE41_out1),
     .PE_out2(PE41_out2),
     .PE_out3(PE41_out3)
       );

PE PE42(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE41_out2),
     .PE_in1(PE32_out3),
     .PE_in2(PE43_out0),
     .PE_in3(PE52_out1),

     .PE_out0(PE42_out0),
     .PE_out1(PE42_out1),
     .PE_out2(PE42_out2),
     .PE_out3(PE42_out3)
       );

PE PE43(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE42_out2),
     .PE_in1(PE33_out3),
     .PE_in2(PE44_out0),
     .PE_in3(PE53_out1),

     .PE_out0(PE43_out0),
     .PE_out1(PE43_out1),
     .PE_out2(PE43_out2),
     .PE_out3(PE43_out3)
       );

PE PE44(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE43_out2),
     .PE_in1(PE34_out3),
     .PE_in2(PE45_out0),
     .PE_in3(PE54_out1),

     .PE_out0(PE44_out0),
     .PE_out1(PE44_out1),
     .PE_out2(PE44_out2),
     .PE_out3(PE44_out3)
       );

PE PE45(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE44_out2),
     .PE_in1(PE35_out3),
     .PE_in2(PE46_out0),
     .PE_in3(PE55_out1),

     .PE_out0(PE45_out0),
     .PE_out1(PE45_out1),
     .PE_out2(PE45_out2),
     .PE_out3(PE45_out3)
       );

PE PE46(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE45_out2),
     .PE_in1(PE36_out3),
     .PE_in2(PE47_out0),
     .PE_in3(PE56_out1),

     .PE_out0(PE46_out0),
     .PE_out1(PE46_out1),
     .PE_out2(PE46_out2),
     .PE_out3(PE46_out3)
       );

PE PE47(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE46_out2),
     .PE_in1(PE37_out3),
     .PE_in2(PE48_out0),
     .PE_in3(PE57_out1),

     .PE_out0(PE47_out0),
     .PE_out1(PE47_out1),
     .PE_out2(PE47_out2),
     .PE_out3(PE47_out3)
       );

PE PE48(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE47_out2),
     .PE_in1(PE38_out3),
     .PE_in2(PE49_out0),
     .PE_in3(PE58_out1),

     .PE_out0(PE48_out0),
     .PE_out1(PE48_out1),
     .PE_out2(PE48_out2),
     .PE_out3(PE48_out3)
       );

PE PE49(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE48_out2),
     .PE_in1(PE39_out3),
     .PE_in2(PE40_out0),
     .PE_in3(PE59_out1),

     .PE_out0(PE49_out0),
     .PE_out1(PE49_out1),
     .PE_out2(PE49_out2),
     .PE_out3(PE49_out3)
       );


PE PE50(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE59_out2),
     .PE_in1(PE40_out3),
     .PE_in2(PE51_out0),
     .PE_in3(PE60_out1),

     .PE_out0(PE50_out0),
     .PE_out1(PE50_out1),
     .PE_out2(PE50_out2),
     .PE_out3(PE50_out3)
       );

PE PE51(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE50_out2),
     .PE_in1(PE41_out3),
     .PE_in2(PE52_out0),
     .PE_in3(PE61_out1),

     .PE_out0(PE51_out0),
     .PE_out1(PE51_out1),
     .PE_out2(PE51_out2),
     .PE_out3(PE51_out3)
       );

PE PE52(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE51_out2),
     .PE_in1(PE42_out3),
     .PE_in2(PE53_out0),
     .PE_in3(PE62_out1),

     .PE_out0(PE52_out0),
     .PE_out1(PE52_out1),
     .PE_out2(PE52_out2),
     .PE_out3(PE52_out3)
       );

PE PE53(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE52_out2),
     .PE_in1(PE43_out3),
     .PE_in2(PE54_out0),
     .PE_in3(PE63_out1),

     .PE_out0(PE53_out0),
     .PE_out1(PE53_out1),
     .PE_out2(PE53_out2),
     .PE_out3(PE53_out3)
       );

PE PE54(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE53_out2),
     .PE_in1(PE44_out3),
     .PE_in2(PE55_out0),
     .PE_in3(PE64_out1),

     .PE_out0(PE54_out0),
     .PE_out1(PE54_out1),
     .PE_out2(PE54_out2),
     .PE_out3(PE54_out3)
       );

PE PE55(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE54_out2),
     .PE_in1(PE45_out3),
     .PE_in2(PE56_out0),
     .PE_in3(PE65_out1),

     .PE_out0(PE55_out0),
     .PE_out1(PE55_out1),
     .PE_out2(PE55_out2),
     .PE_out3(PE55_out3)
       );

PE PE56(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE55_out2),
     .PE_in1(PE46_out3),
     .PE_in2(PE57_out0),
     .PE_in3(PE66_out1),

     .PE_out0(PE56_out0),
     .PE_out1(PE56_out1),
     .PE_out2(PE56_out2),
     .PE_out3(PE56_out3)
       );

PE PE57(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE56_out2),
     .PE_in1(PE47_out3),
     .PE_in2(PE58_out0),
     .PE_in3(PE67_out1),

     .PE_out0(PE57_out0),
     .PE_out1(PE57_out1),
     .PE_out2(PE57_out2),
     .PE_out3(PE57_out3)
       );

PE PE58(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE57_out2),
     .PE_in1(PE48_out3),
     .PE_in2(PE59_out0),
     .PE_in3(PE68_out1),

     .PE_out0(PE58_out0),
     .PE_out1(PE58_out1),
     .PE_out2(PE58_out2),
     .PE_out3(PE58_out3)
       );

PE PE59(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE58_out2),
     .PE_in1(PE49_out3),
     .PE_in2(PE50_out0),
     .PE_in3(PE69_out1),

     .PE_out0(PE59_out0),
     .PE_out1(PE59_out1),
     .PE_out2(PE59_out2),
     .PE_out3(PE59_out3)
       );


PE PE60(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE69_out2),
     .PE_in1(PE50_out3),
     .PE_in2(PE61_out0),
     .PE_in3(PE70_out1),

     .PE_out0(PE60_out0),
     .PE_out1(PE60_out1),
     .PE_out2(PE60_out2),
     .PE_out3(PE60_out3)
       );

PE PE61(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE60_out2),
     .PE_in1(PE51_out3),
     .PE_in2(PE62_out0),
     .PE_in3(PE71_out1),

     .PE_out0(PE61_out0),
     .PE_out1(PE61_out1),
     .PE_out2(PE61_out2),
     .PE_out3(PE61_out3)
       );

PE PE62(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE61_out2),
     .PE_in1(PE52_out3),
     .PE_in2(PE63_out0),
     .PE_in3(PE72_out1),

     .PE_out0(PE62_out0),
     .PE_out1(PE62_out1),
     .PE_out2(PE62_out2),
     .PE_out3(PE62_out3)
       );

PE PE63(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE62_out2),
     .PE_in1(PE53_out3),
     .PE_in2(PE64_out0),
     .PE_in3(PE73_out1),

     .PE_out0(PE63_out0),
     .PE_out1(PE63_out1),
     .PE_out2(PE63_out2),
     .PE_out3(PE63_out3)
       );

PE PE64(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE63_out2),
     .PE_in1(PE54_out3),
     .PE_in2(PE65_out0),
     .PE_in3(PE74_out1),

     .PE_out0(PE64_out0),
     .PE_out1(PE64_out1),
     .PE_out2(PE64_out2),
     .PE_out3(PE64_out3)
       );

PE PE65(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE64_out2),
     .PE_in1(PE55_out3),
     .PE_in2(PE66_out0),
     .PE_in3(PE75_out1),

     .PE_out0(PE65_out0),
     .PE_out1(PE65_out1),
     .PE_out2(PE65_out2),
     .PE_out3(PE65_out3)
       );

PE PE66(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE65_out2),
     .PE_in1(PE56_out3),
     .PE_in2(PE67_out0),
     .PE_in3(PE76_out1),

     .PE_out0(PE66_out0),
     .PE_out1(PE66_out1),
     .PE_out2(PE66_out2),
     .PE_out3(PE66_out3)
       );

PE PE67(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE66_out2),
     .PE_in1(PE57_out3),
     .PE_in2(PE68_out0),
     .PE_in3(PE77_out1),

     .PE_out0(PE67_out0),
     .PE_out1(PE67_out1),
     .PE_out2(PE67_out2),
     .PE_out3(PE67_out3)
       );

PE PE68(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE67_out2),
     .PE_in1(PE58_out3),
     .PE_in2(PE69_out0),
     .PE_in3(PE78_out1),

     .PE_out0(PE68_out0),
     .PE_out1(PE68_out1),
     .PE_out2(PE68_out2),
     .PE_out3(PE68_out3)
       );

PE PE69(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE68_out2),
     .PE_in1(PE59_out3),
     .PE_in2(PE60_out0),
     .PE_in3(PE79_out1),

     .PE_out0(PE69_out0),
     .PE_out1(PE69_out1),
     .PE_out2(PE69_out2),
     .PE_out3(PE69_out3)
       );


PE PE70(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE79_out2),
     .PE_in1(PE60_out3),
     .PE_in2(PE71_out0),
     .PE_in3(PE80_out1),

     .PE_out0(PE70_out0),
     .PE_out1(PE70_out1),
     .PE_out2(PE70_out2),
     .PE_out3(PE70_out3)
       );

PE PE71(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE70_out2),
     .PE_in1(PE61_out3),
     .PE_in2(PE72_out0),
     .PE_in3(PE81_out1),

     .PE_out0(PE71_out0),
     .PE_out1(PE71_out1),
     .PE_out2(PE71_out2),
     .PE_out3(PE71_out3)
       );

PE PE72(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE71_out2),
     .PE_in1(PE62_out3),
     .PE_in2(PE73_out0),
     .PE_in3(PE82_out1),

     .PE_out0(PE72_out0),
     .PE_out1(PE72_out1),
     .PE_out2(PE72_out2),
     .PE_out3(PE72_out3)
       );

PE PE73(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE72_out2),
     .PE_in1(PE63_out3),
     .PE_in2(PE74_out0),
     .PE_in3(PE83_out1),

     .PE_out0(PE73_out0),
     .PE_out1(PE73_out1),
     .PE_out2(PE73_out2),
     .PE_out3(PE73_out3)
       );

PE PE74(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE73_out2),
     .PE_in1(PE64_out3),
     .PE_in2(PE75_out0),
     .PE_in3(PE84_out1),

     .PE_out0(PE74_out0),
     .PE_out1(PE74_out1),
     .PE_out2(PE74_out2),
     .PE_out3(PE74_out3)
       );

PE PE75(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE74_out2),
     .PE_in1(PE65_out3),
     .PE_in2(PE76_out0),
     .PE_in3(PE85_out1),

     .PE_out0(PE75_out0),
     .PE_out1(PE75_out1),
     .PE_out2(PE75_out2),
     .PE_out3(PE75_out3)
       );

PE PE76(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE75_out2),
     .PE_in1(PE66_out3),
     .PE_in2(PE77_out0),
     .PE_in3(PE86_out1),

     .PE_out0(PE76_out0),
     .PE_out1(PE76_out1),
     .PE_out2(PE76_out2),
     .PE_out3(PE76_out3)
       );

PE PE77(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE76_out2),
     .PE_in1(PE67_out3),
     .PE_in2(PE78_out0),
     .PE_in3(PE87_out1),

     .PE_out0(PE77_out0),
     .PE_out1(PE77_out1),
     .PE_out2(PE77_out2),
     .PE_out3(PE77_out3)
       );

PE PE78(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE77_out2),
     .PE_in1(PE68_out3),
     .PE_in2(PE79_out0),
     .PE_in3(PE88_out1),

     .PE_out0(PE78_out0),
     .PE_out1(PE78_out1),
     .PE_out2(PE78_out2),
     .PE_out3(PE78_out3)
       );

PE PE79(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE78_out2),
     .PE_in1(PE69_out3),
     .PE_in2(PE70_out0),
     .PE_in3(PE89_out1),

     .PE_out0(PE79_out0),
     .PE_out1(PE79_out1),
     .PE_out2(PE79_out2),
     .PE_out3(PE79_out3)
       );


PE PE80(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE89_out2),
     .PE_in1(PE70_out3),
     .PE_in2(PE81_out0),
     .PE_in3(PE90_out1),

     .PE_out0(PE80_out0),
     .PE_out1(PE80_out1),
     .PE_out2(PE80_out2),
     .PE_out3(PE80_out3)
       );

PE PE81(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE80_out2),
     .PE_in1(PE71_out3),
     .PE_in2(PE82_out0),
     .PE_in3(PE91_out1),

     .PE_out0(PE81_out0),
     .PE_out1(PE81_out1),
     .PE_out2(PE81_out2),
     .PE_out3(PE81_out3)
       );

PE PE82(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE81_out2),
     .PE_in1(PE72_out3),
     .PE_in2(PE83_out0),
     .PE_in3(PE92_out1),

     .PE_out0(PE82_out0),
     .PE_out1(PE82_out1),
     .PE_out2(PE82_out2),
     .PE_out3(PE82_out3)
       );

PE PE83(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE82_out2),
     .PE_in1(PE73_out3),
     .PE_in2(PE84_out0),
     .PE_in3(PE93_out1),

     .PE_out0(PE83_out0),
     .PE_out1(PE83_out1),
     .PE_out2(PE83_out2),
     .PE_out3(PE83_out3)
       );

PE PE84(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE83_out2),
     .PE_in1(PE74_out3),
     .PE_in2(PE85_out0),
     .PE_in3(PE94_out1),

     .PE_out0(PE84_out0),
     .PE_out1(PE84_out1),
     .PE_out2(PE84_out2),
     .PE_out3(PE84_out3)
       );

PE PE85(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE84_out2),
     .PE_in1(PE75_out3),
     .PE_in2(PE86_out0),
     .PE_in3(PE95_out1),

     .PE_out0(PE85_out0),
     .PE_out1(PE85_out1),
     .PE_out2(PE85_out2),
     .PE_out3(PE85_out3)
       );

PE PE86(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE85_out2),
     .PE_in1(PE76_out3),
     .PE_in2(PE87_out0),
     .PE_in3(PE96_out1),

     .PE_out0(PE86_out0),
     .PE_out1(PE86_out1),
     .PE_out2(PE86_out2),
     .PE_out3(PE86_out3)
       );

PE PE87(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE86_out2),
     .PE_in1(PE77_out3),
     .PE_in2(PE88_out0),
     .PE_in3(PE97_out1),

     .PE_out0(PE87_out0),
     .PE_out1(PE87_out1),
     .PE_out2(PE87_out2),
     .PE_out3(PE87_out3)
       );

PE PE88(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE87_out2),
     .PE_in1(PE78_out3),
     .PE_in2(PE89_out0),
     .PE_in3(PE98_out1),

     .PE_out0(PE88_out0),
     .PE_out1(PE88_out1),
     .PE_out2(PE88_out2),
     .PE_out3(PE88_out3)
       );

PE PE89(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE88_out2),
     .PE_in1(PE79_out3),
     .PE_in2(PE80_out0),
     .PE_in3(PE99_out1),

     .PE_out0(PE89_out0),
     .PE_out1(PE89_out1),
     .PE_out2(PE89_out2),
     .PE_out3(PE89_out3)
       );


PE PE90(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE99_out2),
     .PE_in1(PE80_out3),
     .PE_in2(PE91_out0),
     .PE_in3(PE00_out1),

     .PE_out0(PE90_out0),
     .PE_out1(PE90_out1),
     .PE_out2(PE90_out2),
     .PE_out3(PE90_out3)
       );

PE PE91(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE90_out2),
     .PE_in1(PE81_out3),
     .PE_in2(PE92_out0),
     .PE_in3(PE01_out1),

     .PE_out0(PE91_out0),
     .PE_out1(PE91_out1),
     .PE_out2(PE91_out2),
     .PE_out3(PE91_out3)
       );

PE PE92(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE91_out2),
     .PE_in1(PE82_out3),
     .PE_in2(PE93_out0),
     .PE_in3(PE02_out1),

     .PE_out0(PE92_out0),
     .PE_out1(PE92_out1),
     .PE_out2(PE92_out2),
     .PE_out3(PE92_out3)
       );

PE PE93(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE92_out2),
     .PE_in1(PE83_out3),
     .PE_in2(PE94_out0),
     .PE_in3(PE03_out1),

     .PE_out0(PE93_out0),
     .PE_out1(PE93_out1),
     .PE_out2(PE93_out2),
     .PE_out3(PE93_out3)
       );

PE PE94(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE93_out2),
     .PE_in1(PE84_out3),
     .PE_in2(PE95_out0),
     .PE_in3(PE04_out1),

     .PE_out0(PE94_out0),
     .PE_out1(PE94_out1),
     .PE_out2(PE94_out2),
     .PE_out3(PE94_out3)
       );

PE PE95(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE94_out2),
     .PE_in1(PE85_out3),
     .PE_in2(PE96_out0),
     .PE_in3(PE05_out1),

     .PE_out0(PE95_out0),
     .PE_out1(PE95_out1),
     .PE_out2(PE95_out2),
     .PE_out3(PE95_out3)
       );

PE PE96(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE95_out2),
     .PE_in1(PE86_out3),
     .PE_in2(PE97_out0),
     .PE_in3(PE06_out1),

     .PE_out0(PE96_out0),
     .PE_out1(PE96_out1),
     .PE_out2(PE96_out2),
     .PE_out3(PE96_out3)
       );

PE PE97(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE96_out2),
     .PE_in1(PE87_out3),
     .PE_in2(PE98_out0),
     .PE_in3(PE07_out1),

     .PE_out0(PE97_out0),
     .PE_out1(PE97_out1),
     .PE_out2(PE97_out2),
     .PE_out3(PE97_out3)
       );

PE PE98(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE97_out2),
     .PE_in1(PE88_out3),
     .PE_in2(PE99_out0),
     .PE_in3(PE08_out1),

     .PE_out0(PE98_out0),
     .PE_out1(PE98_out1),
     .PE_out2(PE98_out2),
     .PE_out3(PE98_out3)
       );

PE PE99(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE98_out2),
     .PE_in1(PE89_out3),
     .PE_in2(PE90_out0),
     .PE_in3(PE09_out1),

     .PE_out0(PE99_out0),
     .PE_out1(PE99_out1),
     .PE_out2(PE99_out2),
     .PE_out3(PE99_out3)
       );



assign data_out0=PE00_out0;
assign data_out1=PE01_out0;
assign data_out2=PE02_out0;
assign data_out3=PE03_out0;

endmodule

