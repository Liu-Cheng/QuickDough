`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IuVM5cUtmUQKgTBX7HKDmAT1YvCAn3gPWTRIcJbentll9fNGh9qKWzclus07vxZbvEZH49G727Hp
K/1Dcy0Gjg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pjFrFtabU6Ur8yA8axpBAS/6vABn0s5Akgw0WazBdmxD71+6StDGi/Bx4QL0BkkNNKkDFrDazxt3
IlNaTnzFw1zqKupSfp4yd1jSKCOFfeu3Qgm8mU7TtVTlYJBt32eKWxkirwexrxwAbEg2XW3T0Jek
Yn27OCdgcKdq94aZ08k=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mFBaaqTk6WujK6m41XGuotXsDplj3ilnvg4jovrY5HWjDlNf4lZI6BludVXW6DRreoxTQg2lx7qP
06IyzAzT6wbFa/rwHEtllH/B0yvuB4ZPW223Zp8AK64j61t7+tOuZX3qCDNRUleGw8KqS0WmUjmz
9a4cz/51klcPgO1miwM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q1x3d5RSu5KDehhgH7qcvqPLNq5cPlzirHId1/D5ljTL1hlPrGSgakTWd4ukrQFWKjS5CA1/gqbN
3w7XBYdSAtEjz7zhcIvAQqj0awdn++yJqRY9r4q77/tWPDo/dsx7Vi/CSjqcM2CpbdHSieE2Rn8t
T+FtAhbxFntvgt4F+XgzXXZWU3Q8NwmgHCnauQaiY9v1Jmh0j+AzrFymmW9bmMaAzylNmXG6qi1p
jrPRltaCAoUrnasCdszukKo+d+LvaCVLm6+diTsVRBT3vogtqBFDCW13sAouxJM+gvWyPxlTHPil
dt4Py1wP2Php8/2AQ0SAKkMskkajvR5QqiLmQw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FoVq1Zhjl4mDZCIqBHcehAw005mVLHybVZ9u4ZLn8BYCi/MhJPxgZecQYmqVZ8YBtv+U8tA3ZcIF
lExV/c+rp+VM2Q/j8GTBVFSz8yagdCv+2hP+jluejIPCxVsMiVIEqDpLsX1liRdbWzP2TmEOf7HB
gLvh6PIpzoSvS7uUPxfxTioSnXhDLzQhki7HRLDLB1SMZu6VdBEVoxcvOAKCZz3jd2rZHEqEFw9m
v3Ir5YbUyDuVxIUBezHIBgUws6aLHk9QRZ0vfrEfQwkaudLAcPGmjRqMf4frVvWPB6ZHEMlSqS3L
Oxmj2TotaCom0jcmktsDLCx6RNuvC63Lmhn4IQ==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
b7aqdpotXnkMc4G/M9sdZ8HR6YofY7osQmQe9KNO0CqX4QxV4I0cZ1/m/dS4Tj5OtH2znt7R5Xrn
DXfQSD/hBpwaA87k8AKlhK/sA9/90l5N32YWIaT0qktjHwSJkNCWsF6N56H3mHWA/O+jPz/GYXmQ
WF6WSWMGZ5nYNw7mnYtCpTUJcdqYLvKhmwLBNnzvoXxfXi2ESD/A5OrxRi4XtQ99o0IRQ3oAU/IM
s0maZLuUWpeLZY2T8f0rGGgEGgjM6WqHeFsRNPfpeaxpTzqOxHz8RHi4t5VaVoLLQaNw9s70xOGb
L+VKDYcq2fsmW532WGSy9hqtkJrubwvPYIOTLQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17440)
`protect data_block
UlqCvAbx8AFHB1yGL7TND4VaREf0uBUpH9y//QX27Sf/ahjF8t20rN5tZhqlzApksuUKAFiXNUCr
TRMuzC/ZdwKX9i+EqQ7WRMq3TPmYaL5B1MmpF0O/RviaK1nKfn/369Gfh+NLprykd5xspTeFiIzi
GtJ/MybhGk0ejWPgEItZjb12PN9b+Pe4Jg7TSenC4NLPh1riG0XC0ZU/TkJTzkHz+elZd8GxFTPm
KBf7RVgkXp1aVyZPaZ7iebpJoCsI7q7GiiEL2+V0DCw7taGIWRwkTvsgnpcfclNaDgMV7YJnuG62
O1Jyuxf3cBl59t882dVJCI+9RpPuW4hN1GcUOUlZFBqin4Iwam9ZAIbBfJXMTvQWFlkeD6dtkj3d
wS/MUA0rOE2AwS2yzj6R6hzLnpIau6evDVD+oAFt09A8C+xGKI/k191lvx/RB3j6yTp6n4QMYPVV
+f/ohCZeG9fEuuUnGW2fdRBxGNX+RBoAHK9QdkHSJXoa1VFSOeqUZNBTEcSBKvzggfZ23qxca6aG
pisQHBf97ObAbeHE8UrNzDo0OxDVEv4j4Bf0fOLKir6MQTjXgIjl6Un5ZcfYRUd916tcxBU5fu+8
nXI9Pd5IZfyxbT8vmmDkygvDLOhPqy/tm4NGbgf0DaCqTqRICXX2AF1+0hioOf+TQMs+kVfQbzb0
DHmY6gcLwMqvvsE5zNMWMZKeg2c+x/ysBIzk6UcLgrG3JqBBaXbBNQQKbEkGUV1ox0SIlR7HkjvC
54itxdSEjisyS3BNVNI1FVO5HAbIydnp3mEtjbkCK57CznC3hLqofv1LpKQw9o09pgG7D7ChRwrd
hFDkPSUerGa49ab82rNxYqRbqpUwWL6sUlgXdYvD+a5MbOxmOfUHdFXWt2Xu4uJOH8MySJcfusLV
8VnEt6bSDbPQExQAtfLPY/1qzDqS+ZLT0B4zWbTudwME0sneKTpZwoli0O0jQ1HF9f1B6OJPL7UK
r4/8XI9365zgS65q6UXLlDi1frRsArTnNBtNyDalhHyEB4P8EIWFwbv5wbXaKARJXoYmD8RlQizp
TraOiwA+Rd4cRw3Ma4xiZYQFsdns6ZauZZwxvR595l2hhICGeH2iViRypTX66g9fN2l1jhTAPCY/
/yLIZ69uEcJiYlJt6+Hmsbb4vHwEF8vWxEPdKEwLAEB9aR55L4uB/NZRAGHQqwXOeNXzuihoVSxg
ptGuF8snUIHt8heyl5t4O/QpXykENk+yY3T5Anga8WuRl4+mtTBg05W70p7+jJYI56UmUy3uCrpE
wBDTNRgctXK/rIZMZQKRedMgM5s7/oojmP6S5SMeMgjn2fqTv/21Taqf6ZidjCcI9X38TIYj+xE4
yN6RX57zPCvd0uI8JWgYX/u8CNSKKPs4QIVccBV7Uagf2fMRPy3m3dwRksHqVR4Dbl0pDf3v46Fl
1RKNyQ0Gh4Nzhu/6WLg0Z4MPknLx2QXCbFprv/KTp315pRgmDvN4qaT/vIjK+Huf8UDT/HKTpoIa
RodkfErSpmLNtbk1nZqvhlvFy5dSuCeq/3Xf77wZ3jSx8X10zeEsSz5QBp5UvyKzD9vqOUZIpmic
ozNJmpkRZcN/bWecQioGsQbYkkXd8+UYVzRz5uc6ajoFpN2aT/dAHKedfGAoF0jJuYmyEikzQ45v
hw64JBnKOTTa6xkW5zt5WnRecP/egWwo/yPxeU0YL2tU6ipWtuxegOVRJEABOQYTwk2snZSOcJ3Z
DmiYg3ECnomBW68TMfr5p4Eg5vtp2kryfjSwrA37WXP+CyQl53LFznSSwnN4m/TcJHc4RN8kViiu
9/5iUvXrYUihmfIDzmLGPf3Kt9iaVXDZvNTq+vV9oL5KNHdRMm7maMJIdL8pBA+8yssrN/VcpQe7
D075cvW5lHVnceFI84ixG5Zg3u23DLDiM1u+UfA6Z2VE59BYQD0ts74Eqj2cIvwEmbAosL0ORwVE
pOZaovpfXBubPhzDqBj5Bf+Dg8xy9HA7+bEYF9kKAImLLSCKMlVYwUaHKDd90b214yrdTCA49xA+
oUtNTVicShaGK7V/ir0HPjr6yrLkruJpqul1ZBj2iAFvs9a8Os3JONwEPO541sAiD+tuS3RCCj2z
CJ2M3O20OspvQ6XwbR3xz9cRog/NwovUi+YLQYAiyCsB19s10OgbUbI3qTCVUpNlN86rnNzofDjH
TBvqKrFi+dOA6jKpXq2looHlr1CpHUCP+KwsO/uiKQgUIGyOs4nlnPQNZ05GHxpdeVQ8hpzOeRgT
NZDtrV4nhb72DgoLlXvXn52PEtsAqROc3LJwUGifhR1Mg5jGEToweolnlHSmxDKim7oSkbuYdqZ4
nJpF2irVHUMMGvpikCR2GoI+rYuGrp12nY0thOi7aoRgAhv33DygOzRuXeKN+XpB+4mFfBL59ycu
AOoDruq2R6PGiuJpYAwtWZlUP7mFzZKDvIGr6lQVRPYFxQPQd+uoe+31AS24YJHIi2906GjCt73V
/KMWZKF73z9U10mcQhtRpSTxztGG7wjQa6N/9Ew/E0oSGPHDF6df0WUdfsN7iEsPLdJUswG2dfdF
1gOhK+Uv9m4r97zQSGI9I9iJyK4k/80CWnjjBGHIVR0kxQohM5NAQsZ0H+39Ti7RzhWYj+qJ5WXe
w+UhllIoPmJm2lIvKUBLb8QLiZhd5/u8VOCHlzg9qQOAw6mYVEBRWSu9tHjzCzhjwGwhFINpkTln
mEgbjhGYSdR3qMUuIb0AOU+pKSWglLpDq8wv0Pfdr1H01tkqV0NHmtAsWFw3n6GcsGqpZeH8yozP
1yFcFhvVJsbfuXNsAS2uEemMX7miesx/LDeZhTvURyHhiVNK+GuLLkRVUL2tp4nkGs9UGQDS9ca5
YnJHjBX0vnNr2xK+avf/C0+1+IPahn0l0LDMgIBugJAN7CPxfMWmNIG2BJadVxK+lEuqYhiPj2FU
iEDsnM9ch9f7puwID9flJRrSvii37k31f9AVzcY2UkoQd80Bg5LW7DJuC01yKrvr3mxGK9t3u1fn
RM9JcDiHFV7MKXiajcXiuG4wvlMREPDYKOiuVVsuEhstAMn0TRLxQkz4iwcU9ykai8jq9ZGupqN9
sH9pMkNqwCjjHb6fLWfRHzm2At/hhGWwZ1DwGh4PSMDHJxKKeCGNitZPtx4pBMj5OL2RMy62RvZI
Ti150QW0pYD6KGMwLfRyymv0MVP3GnWEYiskwBA6xxcCc4Dyl1xMwuqGfE/Qehugg2CKN6jQETzz
vOOXtMXmgD+WvvUtv3WqDYunS68exb6qFdl/g8IxALENF+vgnzB2reLy2xfxVdod5nO5M0mKoLhG
yyuqBQBvgIJnWoPPuX5SJgO39U+TiqiHvSbAMIowCsF1G3X9bi2Jb4yzlEE+LFCSBZteimeYPf7j
TpQMxUGYJIPR/WyX+9lGnJbonw6tnb+Tzf+B48JugFu1Tl2AVoYiGrH7l/y3wRexSTumHN5Ci+rm
eqI9BufSj1rHnlh8FFYDpv1LjZMP+zwJyF2lspFi4Bw96cejw0vlfkCOZLdEOJKfngdp5nAxLl7e
oII10KwFGk0C1jkoHq03pRjzLHpD386HN8lmaWH5n5LVtsGpZfVeRAjFoTI/cY8Z5kCzCYR7W3cA
Jg1bV05jDBdRlAV5FBZKkchBZ9OHheuir6p5ih6ZEFiFKqo7L9HgW2hvtJtyOYFXx3A4ON5NMJyW
hZ+d3FxNfQX56L5WF7SNy8wOB4Q4aZnE/SYBOvzWywY9eYPpwC71XvkH7Gqv/yyWWyTzhPZAIR37
JaeAs+VHaSs5oosqKWlQSIaf/D51cKia3y4rGRAfAc61CnUfEqur28aiv4PyJMUyMGdhdkE8WGkE
6mvfsbpzYtkfFj29duO05/SnyN6sWPMmP2rt5H6R/7ZZh5gN2B7ZUdv08TglZFtTk9eoQqeftEWX
KORULzCFfBuBjK2wKgmvoTYsCGK4hdBGvUNMjmNlnB1mAk3xscdyb0m1wxdPCSV1Hpcla/s1Kbkf
XQgGeoRDI7gaOdiENXe8ObJ/1LID4ZKQigbU36u40xO5RmnJ2778eFnJkMr3lUD14pjh63kWQutT
egkxBB4MOqxD79oGHS+uLrr/CuLGMBfIx7ebQHyGVAx8LQTPfUrY8HbFR6GSG/+Fke7u1JTgKPE6
VPNa3f4yymjAiyRIBcxsqSpAlwOyRov2eufROvZ036uSCGPhfbU9mS6Rq1Tri/86lpY6WMnA1wXa
LZH7ngbKfyFv1MAJe1xH5W5sFIL+G7jp8qidPMyBh+OVyFOedR1RAv63pyjnQXeUEXK09PaHFl1C
1MbepDfZE7UIPvoETjVg62qw5+vCqfC6CeQYYmQbVlaKXZuP8Jrpgt8JdtHRAlFq7Bd+C6BP0gxa
WWPlErcmlxLkemCa6TR9K5sQE8Xi+JXDaA7vb0bgn4piBoWMG70cpvlYNY1+OcSmJqHOuNFuBfQ4
kcBk3UeDICKowFftwE80Jlr474SZqExG4d8lXWF0UwlExhmkhIhaJk9PYmsuC69HRrTc6MniiZf9
p4ICgewFI18jH6mVOkCap+tB55lsdrD9+C1f6h0acEhH6ZYM+I4ishMf5FTC4n6TQ82E3nfWAU0D
bC2MzCDaLadsk9NPip6Bw/eb/rC8b2QW52V+NfSxWaY3y4am6KYoYGatq4rodOtAf04GatOzsZD5
ESBPLMvdopljsUVdvHgQNDmhauB62BwM5ng8RiDwTbYIy024JaypVFMrjweHqlOlM25uncVcihvb
9pOt6P1+JW8GzXxDFYbL6C6aZTEAp1BgaWicP9YojbLcjXfwzTRxTE5hB4OOTzRGb4RPWbLFPPgo
0SBp0xqxfrohIFjpREUTe/AZIIe0R19+K6n5LIdkRlQwPLHFqVrvNcgdvmw1CtlCYW5ni3ShOtSs
zzHEK3Fkuf5heb+wxzlhI2YmFZC/f5oCI2gealrlCtEbxCnoE6mg2LwFp32Mh6Tb31jeowXZ0mzG
HD8c9iOMok7aKMALB6jUYjgBeRDmiQKrfzLS8FTDn8NzEX6XO7Nd0GnTSSNV3H8FQ7KpwlX1fyuj
nwLqc7XS+OvtP8RaobNuzu7yrKWDBHBYHWnl2LVF76HZMkVdbQwZPZPhC4aHZFhyf/EN3ssZl8wp
zvIR3pgxYgb0Raz/SnLDyHbcUUlI1UEQCHNBLsO8u5UGmYEgiLTFuefAy+HFpAZuXKks1aSmBdG8
zOEpVy6kt/7zloBFA8Rad/g3XK7FOWLuupN6uRfoqoyNEvSRcvp7BNekgGdD71F/qPEJjER22vt2
u7Dy3S8mMGROjizqiHKCXFfSxyYGnFzxSYixjvzRXENpj0rQoB6IA17ttM+g0WoOHo54949t0hxi
zYjwx1os3N+5TJFvHo41PyZM+8zczau163mmXxg9ItfwqWvsU1gXE6NfJdj3fmXnn/oXoyTAPbzB
zrQaw+9gqPYOJp87xyrYHjKeKUodjG74845VX0VCOTFCObkt4jPIl0XtJX12I2t7eYiKTO/YS77/
Tm17fGDiCzCxjWhpQKdt9lrAnH7PySLW+k88S2w8vRQr1+UgljJqDrhom50TIwznLNkH7y5M/YJ+
e/nZPR6Odb8KzS6l423qAzfEa/3nuEzy5I57/D+VW6ZuZiZWv1i7aCMnxcYnU4C+0OYgdfeBF5kZ
6nJBGA9sIMC5OSl/AltMGJJq5XnfeVUKTDkehe3Xt5H7MUd2ffD6LchpBpCS9eVnktR8cnFnWbcm
ELI8OlS6d8maBMbQXhjGwt2WqTDtnkt2ncnFtrIrsyLWLJWOpiqugxqRl21YrSHGd44L+RfZrT4h
AZRpurYnxA8wzBPrtnaYMEcVcsIYGu1KRLvLwN2SJN97GjyBreFSQY1tPD9aA4vODtYncVoFG5zW
hkbkw1lg+SXwc62yeA3yfVwLyLpdxWZKUUQxtKEezvIjzxqF3TOU/sMZ1tbB6pb7HW1JLjaz6CrO
buINECwphGP3V8q/IP3a/KQBHXY+VcoF3sC0fjOQxE4XvoD7RIJHwLTH9TGVD8wrByk2YSzvbFcw
c1hDtnDbJUf5ZzLvz9JFlT+cz01AlwNzPJGN/mGNymbAeBE3NoJ4GAV+MUu83OVXd6GsQzMsylkU
j8d5ly9UWuoCm/JJmSSU2FZxkPA9qn10hRwsj6eXlwpq+Nhcoux+nymSckUGmctMs7utfeHAZHAs
a9J8VqnulFKKshHkn4JkmmTUKnVjUnUG/wPgzgLICgngwzNBVhm3cmHzpMSDQn0EeGrwNM4XCiMe
IsfCWGLZlQB8fu+IYZ4so7wMZcrBx7wNgTDQOyxe+X6GK5oBYpiz19PAnO0M7/rdY3Gj99Jsy3Br
Ctjza/TUPeQKlkX5GGVjgReYLCQPA/JIZ0GV0SVZBlht+Ld+E1/jSpnlhRtMnlGKQhj85cHHj6V4
oIvMj8weNYnzuDkHXwR7Qx4wC91bBiddSQrjG78OigKL1YLdpML4Ya0RZQditUns3lRPFd1C/+Sl
OlZgI0afYXPznd59NjYz1luHYAXEwlG5FvkuueVcU+OAnMYzhxnNwL0lfkrLtLolsG4gf+UDxZEw
gB8KGOPC0Xkkzk+0ANo+W2XhuT+3+4qgu4+16vu/QWWH9v4kjaAyUqKNlM1dee7FutqrEoDj4DAY
3z60uwDaGvt6IMDv+uGjBE/Va9tU1snAHB9ZnZRIrjE5CGLvG5gFBT9CANsGImx6VhhhJnq/wPIE
WaenFgVD+6KSctf5cu1pM/9oXYVHZnJUn/zuLXYqBhKwS83hK9LhzLNt+iajTPrAkzjVYcqye68t
OLGUJbusYMBQ/QE9BMXOzn5V7tIxaOj5FfNabX3ZkDSv0tWRDMYVbI12ODBmjwHvwdSqj9RxhRX9
wviVyWEVOKKrGklPiEocJag9c0b55jY/WyU5sCQlmyOIsQGbD5wQaAqmaUF5+L2Y+j2BwwFJrwtE
XPqdWIu4UXwvs2MBL9+rR4HhQoQXYmbiauL3fJBf0W81+RGJS/Tqo4CQOD+ngkBoB4AWVtIT+J5Y
Ap1u6Gmw5Ne/TqlkufCNo/Wkn90+XYk9jTiWlXRAY+jTY0ghVStLkOXU7senF34HJxAnb57BXcCR
9n8pF9jANp91dkveN2yphOnmza8cSad3GZQNnUlHJ21hnPwtVV6Vntubph0f6i9wZ1TaJaz0gpQ3
ngqALYOIkZVOkVb9+/w5Gjx1Kz9muDBLuic9L+sKvlXYldrOdtHsr4WPgnkT5Jd2qqSV1hKqSOdq
1nd5H+I97Gei9+6FaLfDtKHmNb7uV88XSmOn9gN8wCP99OmW8cerW/xuXEgJn/4zhM15wS9Xa3mU
byokcriPmOP7OiKCRsf8gPTlCvFo5BiPGfnd9SfReUCgqa/UE9kJubLnUIAeth2nLLNnHihaJUZJ
qNWoBDW+b3sJtCygSbo1iQQ4EimwgwM7bgfpjMUXaDAMCD/qlpZLg90ylNe040BtUKPPKDSIeZKF
EP5flB0xGqFQ5fyeGWshaTmviJabjM4FLa5HUgD4Vjodzx38tyv2Cwlv72zjR4p8or7jol9Y56SY
MrX6O4Jq7s5kdkqSumVqctglr/IT2RqrTu8ItwVtRDxNJkjoPq85eP0Pv6w0C5OWQCh7IpFPlpc2
IiYrhw+Lu1c9y4xddSYkawBINeD0SUr9MrfiTJubVh2Lqs4jFg1LUEi+NghQyVorOco9s1Cu9MIe
pXw5GUM2vsSPPgNWZAqcW7amSnSFazDFCMpY8FR+RIj9GWEE3XLrB9J413IGzXJgVEfd+s7xes/8
sYIKIkTe9j1veFAUDJoC5fRQwN1Dv7AImZDmrJ9JRyTYZpsdZ/TKKGUTyVmQ/d951Hf9e0VZW+bu
sEdl6ofiS0oMagonziYgkCmoTZ3CH3WBHw6cCM0Nw0bFzaIMvoQCCvtitT0NxitUF9a4Y4Csvh7d
CKnOm5lGKrNK/BJ2YdfOKQ0KH1rw5xALNQ/e9gppHtdUnXLdxGm2/XnvRdRcCHxyXIzlrtG70kCQ
+vpG93EDp+SrJErtrybfscluiiXwDextapPwXEcRygg2U99tEh+A0ubUC3BUCxXlHLp8D/ET1OBY
zSpg6a0yfPIpoJJjkdPZbd1QrIc0RQ0etcx0WmGWkkr1Oo/2NUSYyLiHgCl7wUuulD4vpZfRWW42
Z/5WRCLV5oWcNo20qc88PEupg05hz7PgGZRlnBfQp6iRgzacT4Ueubw0T5PnjcKP4CT9LniUSrpR
cRjHnLb+NqLGgXpXz7MeW3424qtdZGiRh8X4KYLnfY0e1bowj5stJdXEm76DV1tmen2y3809XyEz
Ajme6sikd09VulJeuDHrMfBC27278oL3nPhxQ57ioNY8MjKyRVVwD+ZTkyfQZk1AbsxqjbhydBNW
M/96Pxq2vkCvDa9isQgXKCKsMc1NB/8zwAGo/G05LEZN6eZDpbYPh8notdnn4HBwkywANaDU6ijp
5UiyzqmrCsoxyftFbYOc4fSeAUQgLTIutV2AsuaVDsE3BbFLWHEP57a+OBRPLOQB2DysUhh4jvId
hzjqorqd7Fa6XBdNNgi+vx7/CUGBCV8peFuIKAfy5hfYJU4eTy7MIp0xULLalDbFEUVaU/UI/fDg
B/LpVbj/vAQqfIVcn+WO56YngqVAxe8zhLkUBwjrPJFA+cFHEBBRasBWDIeCc4cJQw70pCRZ44VI
OPPvm5wq0zhvHTGk7sf+rUXwJUdZhtCiB5IfEQaKPD/T5g8+io2+j9r1oz9kJTtpdJpUDJ/Cet1C
HcCJ/xsnmpbpfHAC5qkFeG+mK7RC1+555Q5Gsv/+aL1uBK28tfwfutrmtGcwPZLsD6EbAkzsY7gr
PCJG1ET4UTPXl/3fFCXolNqXbyjz0IEKFuspcsWPPMC27HaeaBPwwhCmzQSBmYH+C3WjE4BLnVpi
h2qNGnQL6Hl78rcIHmboNCmrQti2qVt1xT7PBfJjsURbaRZNk0IPB/KNsVBUDDfNM9HvCL8ybPXu
carEoXXrl14OKRfyxIB/UK05S+10J8uuz9HoFRzho6Ttee1jbVe1ht7mLdCjY2+uRVdHX3f5m9aK
dZYVzb1owAdXganwp7qLbKWBg6FoFSUSVM+tK50kmfXrOQXYod2xHirrWoos8TC0/0+hh8ksNGKF
vrQ375uKNov6hO7eh5jZPlicVqAOYCMGGwhYEEWfcmOtbNaOJ6WD5ErXW+N9DJt2ysJnXraMYros
kyNF8XUdn/gBCl5mqpbaAkm8ZPG/iSR+xk/bww+zuncGjtpjAl89mwxwRAj2KcVo8JLTvuaHQgWc
fM1ggia3NARYuyo4Vy/Vtqpns2XH9DZRgRyDHeDPXYWgokJM2WU6Kh1ET0xe+gDifu5YhvLa5j17
vMT9wmtlxNoFWEO/yd8gjlQQ4SfyvdueKjcVYqp4MyID7QW5lxvbF534BZcr/BtaxBmuUABD0UPu
VIueJtLDt2y+IVd7vcfEv636Oqk+QwM+kZJuO/MUiiPdGFhDewE6J+UjDOiWjs8T2PXE8PfBKAaV
DDZ/XaEw6+otudXpnJAug0baakyBBxdTrles07UQ7e+nXgqoRkg3T7jz3xyVjfyqiDCAshj5sPS8
My7JhZn4Ud4p2yUFIHazwg2VIuNW42GSKnzWzEB3cZ0/uyQgElmLd2uMuGcmLKo2v8aqPH0NVFIh
z1KqgI5H5i3+S3fPixRqXwFDbcqasTYPuk0r+p4TdFYC2SspA4JiJtEnzvmSTCLLO1TKwSrGBJL5
BGmLCjr7sCcuNDtFNz/QAjZUBGGu4B0muXFpp9r9juTfvEF5nVGuoiu0qHZ36pu/BL5tGcWYEenY
YgfyvGQVhI7kqZ+Td5ggHOsCgMk4MRYtpEPNiCVsIKxLYAu4PT5HuVntImLiVE7evQeRbcisrmfN
k2YBvYPJi+lfqSBSW5pvD+tN7EDTqLEcvNTzt1sJktjz1di/v9aJxd/Ps6CK+UNyv3os4GX5KYYf
k0vm2axG3tcpF7rvkaRYkLNLx5El+6PkvXiFwipu0sSBXR/JXcDJId1O2m0OhIbHWUWXj801arCq
CxaFJfCFQh5ZGIqK5phtFuBhVddnmjh7Lvw4Wwr1Kb7tg2FIN9Ax2/qp28tW7DS2m7Ga89rSKIfZ
98qV4aCwZBGhfYxVsjRCfVIqaNtNrtm6ajWACRj7ETInVul22YM1jAlKxkz5+Gvd/E6hP+KqiPcj
2LV87tWSrMWKd9/jJ7njn9pwMcnzqSq9bDdCYmMxcnXegxsA1xRoXhp30jX2D10EXB4FL7g+Nr7p
VptFSrD5QjnJGLNsYu1VPwjdkmCVre33p+ujSwxzX8mJTTAOEU15/tW4z6cPZrUU3Lsc0GUW8RF9
unWKYwd1QK+wdfIrBCAzxvdVDQA5N0JvMpbGX9WrEnPTeL4iSkTQ+3/NgJcopcpQcOSIZrQ0NW7e
Ggmn0seb4mbjZrnyJLq+lvXHV2NCLMcuvFWwkhRj43/TRW94jFdGVUJzFykRkqp0pzDNkHsCT48b
BoMhjgo/Zk00G1G92E3S/poP1MzalLdJCsXSlUXKXbdVEulznbrQcjWMfijsocYRzyKDl6BAv/GV
vNi0BbpNIQrJ9wAdx3A0Kba/y4lVFCidk5a3V86WwYC3k9nNS0pTxQUNYWl4W9heKaPN8U+z8KOT
sy8DWnRgoqqbTxiDxEdKwB15A7pXyapDcGcuJFu/2F3A9AlmARus1R5PwRRD/WZq2FyOhWjp6bH0
G+sWyw0K5lvG9iti4TXhVSmuLGJy8UssS2iJHFkhnJKSmvu/OxCF1Qso8DG+E2PaKvZz1oSD/3Lb
0zXxJbTNTfGopCZ7tFTppz/SCkRqpMKUJRmwYMy+YGCGTs3Hig/R8+wKEgyvce8tnONLtAQ/YnsR
zV6texSyqI422fo7fussLldrkjrH+t1j9Y7iXW0lWweHlyMVFEWTU8pmGH0WYDxR9Hx4UW5lvwxh
pk2owG0pXsPOY1U0O6uld6d1rIIsxCDQcgE6nX4hr7Y+uYE5o0lRKt6uu1gXO6Srq31Yqr3s30K3
RV4SWPUyV1BHzN1JvX7eReQtAcPmebnY+FAMHHlWRYiU95UqGArB7CCHm+vaChgLMgmTQg6PGtZf
UFcDSz3QwMBJHWDjF4qFLT57ho1yoV99MEvpCscyMhaMYOSPD8d4ziiRXf1X39rpQPwZ0Qur4m1Y
JgQ5KWlp7dbd3Qr2U2OMrOeUAM9p3p9QaK0NvHIUBwm1fSEXzEoxgNooUytPwwL9lRr7gn+/BKk5
hKC0SRaKGXEOUAS2EXKgv1vKoscoBP7yek4Oc0Ae5QqQzCh2uucFTCOYuE5zys6Z7D4Tucau+UIW
KQgPyyqlpYr22uF6YA1YQ7ZK0CJgZi36pmjbt2SNZuW3i/QIHU24DpBkeoAinwPdtthPfxD9kM08
9m/g07LyypqnP6qt7onjn8+ZopA+g2cbpFIQlH72E3fCYjjF9+56A3NCVU3w0sDn2MMnSp66ukUZ
q23e+gDm294RBZAGMZOaNkGtbQvmZEaaoKVoPthOOpH/Bpi+uidNGJ7a2jsousN7a9unq1at1cHn
4uLkJ7onlqhNSTEpGwmJOfxifrE9eRRyBsvBKFHSTxJgCqj3mYURg1cLfNYpeEOcYC28uFG16a2a
LFbUQDlIUGNHYIneuVuJlx30R3VQ/lo+oQoz7FjKq/xoa8lf3hCOr6IUvm62h0KHtMCyCsMgMPq3
ylr6zUarNwo0s10wZ/s2B+uF//gFm4IeW2/3nzF9u0h+/IuayBc0xQyXpwV0Qe+UDxXxUINeZdpM
/sas34gRyng8koC+kmwxyApXPF3xIlcsxk10XspJlI1T0FR96/06lw6308dnro1ezk2TRSI7FwJp
yDZ8xzhYyijunqYo6yQ0ESgG6OVGL7wYoHxznpdi9KCrI9Q4HfBGZtF80zk7DyUk0CIvu/yFuAbC
xbMwK1phrYxfOxVddFQVAPHvLLSJd0w/M5WP6d1c+ixDI7EapgVfFzPvxCgGqyMT+t8Ad+pkh++7
LANIOzCiNYEw/nwq1sFWeYJdtDK7hwWAz2FJ9kSqnuNjToU7o5yeaatA775tZDFzV/Fitfi0fARr
2BOCuSv+0KohZbfu3OHZIntlJuvMzPaL6plDkmjXEp9XMY0XHNq399S6H1IlrVkGZ3utEpfq71F+
ZWyyssBI+YlD+i4kshck3Ti4eXt5UOlfS/zMPox9rTHkl7zWskyH/eyHDeNK9WZSmXI7kBMMOOYL
fmsi2dUmY5UbrW0KqgC4gIW+m3Y+uRKdf8oeY8aDzS2uCMPrgvP5pQkWju5/FKvs9ZcnfBjnzK9/
RgXy3n/8aLcajBWKh6DH7NMdbsh8jyGEVk05PA59ZfGBkzKZuZ2e83xSOjMcDKcCUiC7CKG9coPD
50FdffNGpkml/xvK16MGyw7D1ai8EQx3XPaHIv4Kt0z2RKgW+XN/chUGbnvShH+T6zzCm0BK8Lur
Z4CeVkX5syRQNKj+a/3cCyd93e/7eRYvZSoxSLVRnrrWHcLqcZm5KR09HzLVQeWQ4mGARSRpt3jn
TdXZn5KRP0vchL6TlMdEfG835EpeH8mHvRr6iQLiHs2AbYwOgSe7azvRB6QOHuQinHvcq+UVPvyj
N1NHrQ8JX/cnG8GXWaXmTtlvAVKOXuxk4JvHe61kKlOpzws+zTO94bATuilqEf5UbSMW0/1poVYf
j7xh7+dOmYKW3bJgt/N7rQrSvRH0QR1ebNVHwzAjavJWdJJEL4e7XtGGLLFgD6TN4m4Id5tStWKG
5SnnGSdAp4/6xzyOTIWUgHMZbS6rPb52/DOt/UL+DXjbN1vrDGbBNGUq8tb74v5yObLXQ8V0/aPq
t4ePQkm3w3t010vt7La6pApXqtT9VfIcqVgbdhwxvd2ws5fFQKCE1QrwIca32AUGaKiqzcHkPtjm
sqmY85tGKdE427xyNwsJZXoZMtRe9tUD4dy85XxzCxJskNmn/YQerZjXN5TzJefzJ5JJhJ3j+ceZ
AuJs2P1INxfQzuazIiCEPRAadSyzntYGFwvzn56pMgh1uMBYiEKePuTC8KOtMYkpdCAthG2Zr47J
GL5a53gzupPgy16w5iMnXxB6BXJsIVu3VtFNdhimD324PHL9W4bK5di9TWAKuwVWjcxEe+vxOmSX
YxeotLuROTR4HUX/1a1/4pI4QzAIM1N3t+4MACyiALRkYpqWMRyua0rlRZrIGYOPwoexAAmBKvlW
qaXQfq/BPWb3rEWFRzvzJ74X9yV2b8PnRchN5ZUUdTVmg1BS9+T73pDZSz5MCUAsv4fFg5vJiY1F
8yQG3xJZCN7swmZZ7+0IdzZV+Aw3J/lCb4lYvgNpbIELSMbNh11ARFwIi4lHuHtsF5MxcBzzfhb7
sLDfPNMyBsFtPoac1/OPIqCLjjb2JHiPmWCN7LGadKCvnUlHQcs2nDLPmTJvMhO60TZ6KYxwLR9A
+gL5ty8dwcwJXlGuwDWNllAH4cQtx0RFFD/1ZB86JpKc3cuU1vBhmccQJW7n+NmNfG94YQ3Tl54u
cJQqdajOjGdSzS1OaZD3QIYMX7BHdgDwuCR0TEDXIWY1Qbjwz4Zyq2xgWObSXhOA6zWCf/oO/vfK
uGsBbo9FFdixBEz9DH8+KmG21Y7aYZPYMjHu1NpukBlm5jQvK4pT+ZxxtuH0KeHC1sqU5V5qc54w
gTBLiz8YOfXtkjecHqlLy1LJaZ9Af70dVnYMSmsMGgGpsDBoEcPC8obH7zB9dSN/YF74Y3ahd3iw
ausYVxiqbLyCtH/6x+syv65fAbEX/1crM53guyarEBgTGEoQkrUVXfk8VxUaLnibwrpATiFYOg37
BKHCsD/ZyTfWkP9KXNXEPMAmJQ2yfXp0cc7BVAHXfhHNZENHeTmy5byrlkhK4/EWZouK2Tfyh/FG
OwEigFlZE3ua7Qg5eN0aLA2l9ZgFrXVaWXfMSsyzR/Lz++dwjLoA1vnXsyHgHmOEFRkvzdAZmKSN
RasC0u2wNxYQwLvf7cFZRqpR5tb4i2qJIx+XsTEQuog07Rb+YCV4SkvcNHgw8U3TU7Lz/plqmxOy
jy7Z4GDAlVhU42eedMiy1+zoqQWgwt/3aTvZQaUGlq2war9CHtuNeyVJK3n6OPBCBKgtR04m4ywO
xvhtVcn7XNZM2ueKxl9p82jjNhiUk/cyDeSOqRu1kecfAMEra58uxHCdQm7YXPLeKUGfYL4dc1sl
OfB4b25vk7YXRpUW4kKyE6LpwzES0KrG3lo5U4hBmN4QpycHRkyPtDbQmZyOaU+gSVK5ZZNVF9PM
C42t8xjMxonHux9WvKlWGywnL+P5jRe7gOra6+Ya43r1LIaO498RoO5xHtlMHdpgijXPTmmaV069
WS98lRo8Q7zXKP4p4LuFMkzg7ngP2Pz0e5ls3crpxVIIRlZfDIzfigwkPePUE2PaHUnjB9mVU1iG
yd8NS2fPlBZCcdqfNSMMYTElTFJOTYH6HRS9fMoC6b5uBIucEaGFzOjRpmlJwe7esVZlBSDtuXF6
so7bt2SdSqRVI6cdh8XUel61o/rfOG62h78Y5yZyODSukHdwXOfqzjujS5xW7yU+81sc+Dw6CdSG
WUpDKI0ggoqbggTNjzu7KmDYuBA2InShzOg/e376Z6wuaeLyPTs+RL+jvu9ZMKNwYT2LY5uBtmcG
WyolDypaWnyBABUfRG2GXvmdTtuit7/Ob5Y5/Rigbx2UELddg/otcaIqBq5wg66fsEDZz7QzmwAf
bTv6FqbqqBTcrs04Rg982+BsgL8RVIKenSL5t7TsSUfT9nKADPj7r2YQewV62toZhAfDFSKEuuM6
f7oKX8jv2WkVYUtoY3J8Dvj32YwZTi659GeGJTiJWIjRxFGbvKuLkFT4Au6Jpj80UT6wWrcdQMD6
sKlOFjcTk3mfIqIMaEHAeDF0ZI9CB/D5TapsolCj12VIruf4zGALhe3Un8vH+UeUaCeQ2EWFg3yz
+bLTxA8jCIEYcgjXsXUy+1rXT85Y5oTyRyFyycPJrE2jlpMLl3Ho6nuSUjITuR31uDYh6lH4zGdX
Igm3tf7lLtdVtTe3WahZbZY6TeoUZrZEh18pAupC7IndWEEorNvHE6NRYgdpKnc4PaZTC2DCppe1
/r6z6nYRp9gvs6IJGUBgWBVbRzwFQxHKIj1CWJp3IScUiohaa+AJksqG2e4jcD3ztg5AaUoXluFR
TyKQpZ0V++0DuLLmyPa14gh/w4ns8Y3zXFBr1iw3EAdwIQR/HHXgQbCKBaZyek4NyyEI41jWfsng
OZjlOaOsGRzT6a7eLK4vR9dp7d9o+VrSuDhSQ42JZD3fbVByh5Z8JztfXtEp2XkCq/1lqN6ScaQl
cgay2KNFtZ4SCFgskV4snVnvENYh3slplqZq0rUJ/fWbbudWauhieF66t/FLwER9y8McIrQxZkGE
KX+toRXDYZmko1UBtvsKA+gcXAjIO+8D2b7yW+es/9VFYwkLzHfX5JBsPD8Nr3Gk3ve0o++5pNo2
RXB822ayPF5Od0w0k8uqMh0HPF1H6O64uwUXPOZMbUlA5NeSq+dI+jqD7As5aTWxFc5N3vMP02h+
HLg5Pxwyu8+CAzDntznF0bKWW2nhU6PXxmWyFAzsUK6Iy/W77fxIw3hI6nRDiJx0m/FqBG6xC80T
peyuuLivuouZlu1c2yP2dBBrazUuYNlJLu7gLTdHlAY53hr+MItlxGGQU8Z9wqUJOF0yMUrlBQT7
2e+MRr3hnKLlwfDIas/NcjgEmn19rTvE3UYjpllQD1wGGwTgowGthODtkBKknVIDAoKXkarW7cax
szaRJciUGMiOLIrJNDvoC7wjORNK3aN+TW56Z4mmJwL7uNKg8J3cj23p2t2w+Pq9AQK0Ma1uZuUG
bwN1CpnXxRqIsSkvKzM9RiIW8WgxnzAs9awNf88jof0OCnG7zQV+UF4dYZ+JFkKxI69UuzcwL7yh
JDfSPfnNEcsqe+utBClqE26bdD9q06eDacRPmVxcddD69qvSmQW2TtdHIlZmenLZRkp6Jm2N/30o
eCmHmcW/T4qxrBhPq2KEDbIY4gByVyISt4KPX7dP4L98mOP4hGGgS9E1L6NhJWr9qZSq3VY/G4hJ
8JW2B/tfh0swvi6SCBN3rk+qizzsThdAG+Y/Q4PABpwTpNB+YWJYdcGVnPf9athZI+25tIgVojbv
4rsdD8qNqluEWun3LyKXKSdraFj/A46HRRSMpno2X9IXcLAiGp4ROJQ6tVWlYlVqRaFts3ycpkc+
xzQzBvgPv+VtFNHO3vwGKq0EGOvskoinsrnjLrt8esR23GRq76ViHTz3rPhphirLFMYpiPos0Lmu
Y4VA+p/3vw8YK9Di3rCErh6NrZRgAKNEGrCwDrpZDbRPWXOIN699S2seyV7GP4FZXmfctfD/Cb9z
nKl/UN04YOf6Vc5882wCLIdFhX+tcJH2ldxlD6DFTy5t0A/TmOhxMCmFPcOBTGnf8fvrkYX38sOz
+6vZYjLfajBuE1jZ9nRyFn9yYGmQWtEfhWs1s+bmnmm5jGMr9XK2WoY2I0EALm/3Fjigev6CakO3
8xDXKZR7sPL1mdrVMFy/wR3y2AVdAfnptc3AYVJtuh/w/QHA4cDzW5zFaNx/cijKo9nnBWQrMpC7
BaeylE8QxqiTOl6NW3l8KssG5S0trHhgL2JKfvuz41DmiIIe7WOtSn0PAdXH9DZH5XySZnSVl5/u
5P7ExeySmeEewVYQidm96nHb5c4LqMSDD67p3lvCB/99uA1NPqKjc+d1tTczmiy2jcUZQ1Sj0OpU
/ffudzuaUSdhqylOP05IdlT19PxBctM1IdEPa2wHgiaEDSyzgqumnnamrzi+nwvzFtmf/6Oc1Xmn
220mZuDG4mj/yJQzYG4XAqMhoKjAkhVCVEhoJ5mBP/Oq+NVwk6hlpP7UtJURmil/vnb2z8fcCFjn
6OH5rNwgaSpMUSJvwIl7662yam3R/b5ljHkM5O35eubdlxbp/4BHGw9ihrPRSB0E6AB9OIwr4gtf
qmVFgFVntgyLjpFwO4I96anM8nHJ+VgJ4g2X3sX683HOWku6Ye4eVo/XSFInMovZQxGh250fVWhy
FCekl4eJYR4Ovfu5oVt6Fcq2szSnRJSp6byTLuptzFNMKJL1v3rfzxBG1N5jROkw7IRUiZdI1abL
XIM7bLdNVw1kngGBRE1WEE5HO307ZBzID0ag2T106r7H9dQQSylZgjBvIno3OZgDSqbqZ2ivk+MH
aqomoxr1ZIIqTIq7Ob95tlHZ/W4LtFNDzkC85h/YLONr7vW+IgqrFWwXjVoaaQfjlokemP6Awybf
k+vG2zC3FE6boZkOp5LUVE/1WYNLUwPa56eNuHtVkijTR2WI7TR7fWa17ErAfhTddNgjRccxG4oJ
xNQS2a205LW9svA1dXIhYpkXGcuTSwcTtXuIVNdrDxQXPWw40Y3N/paoRXXhQz5I+suF1G5aaSIx
IoaxeAbivKrIA8I/DWhtwafExIOYlt8IwVuFJ9tKY29C8JDC7z58hIKarXVrN/Z5Wg8s/k1GZLgP
mzAknljEt9FH/7/2hkbQ1+YxN6uWpu7TstBQbNh3PsRoPWe6+mtLjfRqzPTFKjypQ0Fqfmf1aR0P
kvci/dJ0rmRv3iKriJfDW8jHwFACJr2hVs4HuNwifH5d6Yd3ELwrSWhtpDWHr+xU51XDyhQXMxdq
ZMELDJqzbxqRpNi0hlUkZ3nKve24RCVN0jElRYoMtlEKxbgYlOF0M95r6a3Y/LFf7FM7/aA0Brk9
BjSIMwAEBeyH3+mvGclxlTHUAGjYxwMcBi2ZE4n/RbGeOu66Y+bo5GsByhFdZ8c7vQUKlcl4xSrI
Qi4yquBNiefeR75l4JzopeDviO0DAFFCFoKU1M4BIAF/TV0LTW06cyStjXbNRfQdWUPj2/hw/Y7P
mH3rpg7tsWxu/6kjY+zW7BqIyxa0wS5VHJWmkDomLu2bpZkCzqtut0ItGVjWJxmW3UpVZ4BtKv/g
QB47+X8UzzAA/XOLxGz3hwDyZeaTnlm/Ph/XXskKBr/IiB1NQ0QGRqVLMFVThJzM/WdXarJAlyA/
R1KojpXFlKBaceNEUGyku7zexsG2dKoyEKhkAHDEytff46GNx5JBdfBMW+HC53cqZUbEGlRT4YFi
UOMOqrwUDHRyaGTCjDupkXmgyZRRrEmxvsgXD/iAQ18XSt5N+/GLkoUmljUNW9yLoFrZf1xDZFME
Tk+Ka7Ry0evCemCnDXi47KtON1+CvW3aZ4gCBO+N9MxJ8ac3F8SB6RsRnJ2DI4RFjIRqdrcAfVs4
GCyajwQzaEFW5xGzn5oI7iuIuwUzDombxCN0COmM3ebpHPhfXgcXaWAl6Qheb5RtQF9Znfmvyb7m
pxGYOjeVDps3I5fZDw7AlrSTUnm+C8YDyjRmCfuNw1FLBg/0CzIo3OrcW+aFmWoEfNlHGYSEo79o
rmg/lW59h4RaCwVjWKe4ngYlaA7zjEYkctRDmSRqO5XSg3y6e3mt/bvTIKVD7D4cTD9gGZlTfrnL
ImBdGu0ljPGVNifaRqQ2MazUdUZv73IUE/wuJaJEi6iY98+8VCKoEplFQYyLPZnpjaedANDUR+oy
9fd2dX/2H6NRYCMs78Saz6d12744nivz+LO2tYXsn/V/ppCS83vVPFGaR6raJ4Jf59LsrsdrOjq3
fDCWGis9KyP7n3YYDGqr4f7TzCdGKnDzfIKwcGnuIiFktqW/Sa7SHHql0njvUws0T7eVkpnMeeoQ
Z0ABYSRCaTy2YJsFZdd7sZb3WGd7BWY+LAXQK55UYP49hu7lNoqp4E+EWzktgjxNT1tbog+xhLOO
KidVUby1Wuwn2Dt8xkSb0wBtulpJTOuYT36457UgROi0lERpkIfavrv38shDVB0fnHisjnqJXfgB
V6awbbRVTnYgJtrOirGasqmUlJUfEYsUMWQRCMrS/izfAebW/S2yYn00AMvhJ9T7EMGl+9keeznA
dDu6yQVXg9NjAzZ+jK5LDhDWmjpcDiS8g9R/MQ6qEqmSO2pctgMY6RQUe2aieRLys1v+Nw9g1b4v
cOMo2H7wirM+OelPHTJY95J/8IWzU7MsXwRt8P0cEeFJkg40pDWj87w8DnjZOrD2NBr1s9mBDR6s
ev9VitQPO7/MQPVeyUkGKMML/F+9kF5qrSlIXU25Iq2LhlVUlsRWMkYpjfw4WRLMNRYTRXCre6za
iAQZiCVsA5TmYLYvg9LFlZ8nR44u36ICgu5QIaPltkVlwZRCEBLl/L2b8Bgi0g6i3tZfEv0zQP9j
fp+5IPylRCejVYLC1DxyhboEDr9/2NbemTZidvjHtps4WvVZ6c1DIojPyAhnIvcNSiJRwK0C8S6W
AcLjNYeauJ31+ockS4gSXNaokUCM1fLCqwS1KuplmfBxqwfP5JbxTFXRAhg7WG1Hk8IXzjx4/96g
ChSbNnTGKl3SHpwbtX7A4sBmz8hqe5Iqp/5goZayZtwFxyarNBFTzj1KFPIAuOpAjw9yyd3Bp5bo
q20fVV2kC5EBfUOi4csK7BwDSoZOGMADNCVYRhyWgY4NbM3wRzLhC3gFubSjGpb/jkEcCn002131
VMQ8WjeLg9w7k/4B67ibZ66WhY41ptYKsXN7EHGv6jtxZMh4LLJiXD7h20gadtlZxxSzcQLe9BrU
OR579a7bKClB4cx+yxQdkMKBepT3Z85WtX9qjZ5onAEbXRdcrPQEdcBOm3jztxznBFYywXghylPA
FTPEt7r5KjW3Ckic/DORCKe7e0BrRDTbmzqQr46aYg/YBq2eMadxrjDOjm6nV81PN7nCClQUo123
wUBKx6LVBKTeW3leDd3KyImI4sPzyZLd67T57SR7YShMjfhEBXmtnkpohlc30xx4IawTFK/mxCVy
b7fSBZz75BMwYcEr7BE2BiUaEw7/O+05dp93bqTY1eE/+re8Lpio9zKP5cxWr4gG00oPvxzvWQ8w
h7gvInajEn74B7DnSJQfpsed9QbYkJrKPW0jlk3TERy4tZ6Mzv0kDPiai36xVMDW2p0/TUiZT68i
kH3as7/x7IfYL70DOQ79+OJGTI1qAqMjHJ7Ldxmoezpn1/RPIPX+d+RDRQuAaEzy4gUUM38DZTzu
bLAQu77O++wmzc7Lp4wOEAoOpVaymUiIIRmLnip/DP2rJbXrbbCfGhnvfq2AxFfFANrB9paHARqz
RTDP+1ogSU1dcB3ATeIM68AELTP1uzp0++/Kr9tnbuvOdkFw+2iaQJtY/ktdDca5dG+8Pe8jgzV0
YukdtNq2AcfHuRXVJsozkjIw6ZGmfBe4bzYqGxI+vGfk2Om1DjZyVPldvEXac9nDXUWYwwXLSLuj
9EPBK7lT9i75/P3jearRQcvD14zNGAVt1h868DGQeHSd1E07ZAJQ6ABlRsZzUBNKkMhPfHFZ6PHY
y876ey6LMUtYH+mMlOT1ujCPDoPyoQrJZte+Lfofx/AEJ+kGvSH15xr7OEZnw5Hb1DmpUmpZ7yMh
UVxkX7WHXI2tfS3Flo4ZzUUNZrc/Cv98V3y3czgScaQomW5BevVOwo1+LL9N1bXdpv+9zcJc7ldN
0AWtjI/gxpZmeDTqdkXcwE8R8cElD84ib+T1HN/vQmIzkrd4V7fjzHN0ZtycJ5aD/n7IkiUK24OB
lmONm06jt2b0FKLivc1IpWZ7x9er09I+A9oVaZZZUU1ZySnziShWZaTfVTT+9bOwan7rbrxDP/h5
kd1Xrsu3/MvQll9qQNQ4VVweUEDpjondZ4fj2zqSudDDICIQfWLHwe0HAUDaOPMRGFrRwyMsXCmq
MVEWM5p1mKJxdrzjOPPJdoGV1g0lt6egAvS76RzzYkJcs0hkShAAMR3lxh0f1hUSQPa8cyMwyqxB
OLLUinwR5/6aKumUh47RnRrHc7Z2uj+in51aiQ/eX4CJijiRJjD6je6TPnilMRe9oEv58gorFehA
QPfi5grATWrfVgEpYraaRdOUOaW+Ei8PFUeYZVWvkyAvPxonwoVJKcR2pHKWZirj7v3uuMcLNI8Y
/He7MzLQBGbos/S6gAb8JlrzmLTEqPv8zpNGU1Z0PMT8S/2h5Z2yCUbe9feoA3GYJ4jd5YGipG3j
uuKEAvqd+rrxQ99spj4RFy2OahQqLg/YiuOl7X7oB8baNE7t+PgMgYWpokT9cOQP750dpXIpywPR
qqg84HpGRXCD/IddiAyKU3vLmCgEkrudLEKq/drnxpFaPJFYOuvJn5KNtF49E7Q/4OSk7fJSowG1
ltK0M6wSreoVS70Y8lZ4xuTRFoxK4ootX8sVkilrcZ0IwkPodFUQtZvwCl5KTlwtty38bzagG7QS
/930FwSQA8Sb99kOk+20kz8/chZHYOE9QPfckj8oU8s09NYMIXgYwpnucvbJKnruPPd9I4iHcISs
OuLi65DXRwaMOeS9uVYsE8dhoEapC4m0KuDyGOhhQUvwBhGAr2idzXRQStHt8Q2zOsACRbUlmTjM
Xmrrp8u/A1XDaum2weFMwAgHW97drpofJlXiF/3xN4j6kFBTfa6OvkolCofNkIG+sswYz1vMxf5K
CVy+XrdCcmQQMOcYm8QWkxg2xvAi3JBZbsSEJKuAZOYlpxigGblMOM6RqLoAaABrQyo7fY38BAAw
nO+6DQcNQX5Hd4QLbd8xLcJrPBrytSQ3e3hFqTfjQPeqFXx4qA+N5RKdLe6s+i04z/XkTmFxF7Pu
KXOVCUXsyn0cHzecYZoIDPfKyJUFtuYiuOn4D/Bo7P21NLjRrvZ66MbbRPzwegDSBUD4hObVkod/
qZbFQvI/1RzltPGSGhlgq5sET3/MwpwvamzKgMbNiX38b3vI8FiqVugzltnGlw4MCFWoELfgRnhO
9CIydWCkn0ay9wd9hZZYPeYztTw6xIk4k6itjjKCX+p+v05+P0VIA6sXVaKiGwGAGBb2WDXK0FVm
N/Y+Q+mhJYmnRnQK/XhN9ObyqiuzViMQWyxZr5ZXvxfAuYyV6h3o9DZHWLV8OHzmtho+UZcalIZE
7PWJVtDp0UEhwRB53O/S7HDYtqExTyX9QVvcVnOw+uDijWklNhNt03GikKcynwSs4WHYpAtK/xjS
hbSj3yDZ/mWfecEXYOosa9+xfoakLrxZRqV4r6sJ/ziufEWNX6We2zGR9Bjd6RmbcDxVBUSa8SBr
GyovJAWRz6fUfCPeEZKkYJZLAJSt+SyX1JzjWZZIOp0WTRtHMmPSfj9pdeA4RIfBTBGxJR/6a9Z+
KrfPgB+OvDPk/PoEtpNWj7J8Txlck7C+paqE916UHljNkZQ1SKGVgbjs8ekSAxtSqQPxihOycg8T
Co+3YZrCRkzJOxyFPuyRDle3VF1iExGKrWRsj87hCia26vnO2sOHunrNp640dW17IsehQjhXn26Z
lo0X1V1OgjetdGKqXgG9DdQdzKvuBndFUzZmj9h5e1Jxx55Eisq26Qu/MmJgBo41GS4+hDLhYflK
5jOhzl3fQhoEKSSlgLGOg+mN+dMd9faEijIJd6sleV9+oaDJP2H5MCbCQYEv3KDaQT05NNSHm1Nx
fs5aTTg7p5BVklADa3ZHA78z2dbhQK4EZsDqvrmMJzXN+TgB3IBbK/LiwP08fi8UuOd/f3qaNai3
9Ay4jDpfuNroByrR3WWdwBQUuDL2vEG0TQRm9ASoHcZQKTjcUvnfTENY+oT+JiP674CfN049pz+Q
mI3fzmBiPYiaF7j7VyGuvYdHC1n8SbkdkaKPou+fOJaZQDca87tDTlmzEWD2lraXv8v8H9mH7+dq
xLYcu90EOwUBqd2th8xNWu3esKnGAVK+8IKM8A2C7eWzMmUzK+J2vZh6A5M1RvR18CI2kFoLhmef
PCqMjBgx7kIkyLuxRIDnmxeP6PfSIZRnSwhTZIkbDoOxhPHNVcA6yyO/KvSi9PdkrNp2rLfUkXdS
7y8wVVO9Bp7vqFBzxXm8NK/QMrUZGibAyxKNzPFf4icEjbrA/KK0UrIfvZUmtbzWrbFX9vR78RSr
rvnQmeAz/e+dhXbvceJubsEWyV27CG8cNPcXmyzDtLu54dfghThzKgMidP2GFu9+ivp5gJHVztVc
dMv96OUK++hfCsB33FvvR1MEtCeFG9qTOaPgDmo7cZOSsUANreSFZFQ9NUl7c83DmPTs7g/hKQ==
`protect end_protected
