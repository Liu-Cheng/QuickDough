`timescale 1 ns/1 ps 

module Torus10x9 (

    Clk,
    Resetn,

    Data0_Load,
    Data0_Store,
    Data1_Load,
    Data1_Store,
    PE_Array_Busy
);

parameter DWIDTH=32;
parameter SYS_DWIDTH=32;

input                    Clk;
input                    Resetn;

input [SYS_DWIDTH-1:0]   Data0_Load;
input [SYS_DWIDTH-1:0]   Data1_Load;
output [SYS_DWIDTH-1:0]  Data0_Store;
output [SYS_DWIDTH-1:0]  Data1_Store;

input                    PE_Array_Busy;

wire [DWIDTH-1:0]        PE00_Out0;
wire [DWIDTH-1:0]        PE00_Out1;
wire [DWIDTH-1:0]        PE00_Out2;
wire [DWIDTH-1:0]        PE00_Out3;

wire [DWIDTH-1:0]        PE01_Out0;
wire [DWIDTH-1:0]        PE01_Out1;
wire [DWIDTH-1:0]        PE01_Out2;
wire [DWIDTH-1:0]        PE01_Out3;

wire [DWIDTH-1:0]        PE02_Out0;
wire [DWIDTH-1:0]        PE02_Out1;
wire [DWIDTH-1:0]        PE02_Out2;
wire [DWIDTH-1:0]        PE02_Out3;

wire [DWIDTH-1:0]        PE03_Out0;
wire [DWIDTH-1:0]        PE03_Out1;
wire [DWIDTH-1:0]        PE03_Out2;
wire [DWIDTH-1:0]        PE03_Out3;

wire [DWIDTH-1:0]        PE04_Out0;
wire [DWIDTH-1:0]        PE04_Out1;
wire [DWIDTH-1:0]        PE04_Out2;
wire [DWIDTH-1:0]        PE04_Out3;

wire [DWIDTH-1:0]        PE05_Out0;
wire [DWIDTH-1:0]        PE05_Out1;
wire [DWIDTH-1:0]        PE05_Out2;
wire [DWIDTH-1:0]        PE05_Out3;

wire [DWIDTH-1:0]        PE06_Out0;
wire [DWIDTH-1:0]        PE06_Out1;
wire [DWIDTH-1:0]        PE06_Out2;
wire [DWIDTH-1:0]        PE06_Out3;

wire [DWIDTH-1:0]        PE07_Out0;
wire [DWIDTH-1:0]        PE07_Out1;
wire [DWIDTH-1:0]        PE07_Out2;
wire [DWIDTH-1:0]        PE07_Out3;

wire [DWIDTH-1:0]        PE08_Out0;
wire [DWIDTH-1:0]        PE08_Out1;
wire [DWIDTH-1:0]        PE08_Out2;
wire [DWIDTH-1:0]        PE08_Out3;

wire [DWIDTH-1:0]        PE10_Out0;
wire [DWIDTH-1:0]        PE10_Out1;
wire [DWIDTH-1:0]        PE10_Out2;
wire [DWIDTH-1:0]        PE10_Out3;

wire [DWIDTH-1:0]        PE11_Out0;
wire [DWIDTH-1:0]        PE11_Out1;
wire [DWIDTH-1:0]        PE11_Out2;
wire [DWIDTH-1:0]        PE11_Out3;

wire [DWIDTH-1:0]        PE12_Out0;
wire [DWIDTH-1:0]        PE12_Out1;
wire [DWIDTH-1:0]        PE12_Out2;
wire [DWIDTH-1:0]        PE12_Out3;

wire [DWIDTH-1:0]        PE13_Out0;
wire [DWIDTH-1:0]        PE13_Out1;
wire [DWIDTH-1:0]        PE13_Out2;
wire [DWIDTH-1:0]        PE13_Out3;

wire [DWIDTH-1:0]        PE14_Out0;
wire [DWIDTH-1:0]        PE14_Out1;
wire [DWIDTH-1:0]        PE14_Out2;
wire [DWIDTH-1:0]        PE14_Out3;

wire [DWIDTH-1:0]        PE15_Out0;
wire [DWIDTH-1:0]        PE15_Out1;
wire [DWIDTH-1:0]        PE15_Out2;
wire [DWIDTH-1:0]        PE15_Out3;

wire [DWIDTH-1:0]        PE16_Out0;
wire [DWIDTH-1:0]        PE16_Out1;
wire [DWIDTH-1:0]        PE16_Out2;
wire [DWIDTH-1:0]        PE16_Out3;

wire [DWIDTH-1:0]        PE17_Out0;
wire [DWIDTH-1:0]        PE17_Out1;
wire [DWIDTH-1:0]        PE17_Out2;
wire [DWIDTH-1:0]        PE17_Out3;

wire [DWIDTH-1:0]        PE18_Out0;
wire [DWIDTH-1:0]        PE18_Out1;
wire [DWIDTH-1:0]        PE18_Out2;
wire [DWIDTH-1:0]        PE18_Out3;

wire [DWIDTH-1:0]        PE20_Out0;
wire [DWIDTH-1:0]        PE20_Out1;
wire [DWIDTH-1:0]        PE20_Out2;
wire [DWIDTH-1:0]        PE20_Out3;

wire [DWIDTH-1:0]        PE21_Out0;
wire [DWIDTH-1:0]        PE21_Out1;
wire [DWIDTH-1:0]        PE21_Out2;
wire [DWIDTH-1:0]        PE21_Out3;

wire [DWIDTH-1:0]        PE22_Out0;
wire [DWIDTH-1:0]        PE22_Out1;
wire [DWIDTH-1:0]        PE22_Out2;
wire [DWIDTH-1:0]        PE22_Out3;

wire [DWIDTH-1:0]        PE23_Out0;
wire [DWIDTH-1:0]        PE23_Out1;
wire [DWIDTH-1:0]        PE23_Out2;
wire [DWIDTH-1:0]        PE23_Out3;

wire [DWIDTH-1:0]        PE24_Out0;
wire [DWIDTH-1:0]        PE24_Out1;
wire [DWIDTH-1:0]        PE24_Out2;
wire [DWIDTH-1:0]        PE24_Out3;

wire [DWIDTH-1:0]        PE25_Out0;
wire [DWIDTH-1:0]        PE25_Out1;
wire [DWIDTH-1:0]        PE25_Out2;
wire [DWIDTH-1:0]        PE25_Out3;

wire [DWIDTH-1:0]        PE26_Out0;
wire [DWIDTH-1:0]        PE26_Out1;
wire [DWIDTH-1:0]        PE26_Out2;
wire [DWIDTH-1:0]        PE26_Out3;

wire [DWIDTH-1:0]        PE27_Out0;
wire [DWIDTH-1:0]        PE27_Out1;
wire [DWIDTH-1:0]        PE27_Out2;
wire [DWIDTH-1:0]        PE27_Out3;

wire [DWIDTH-1:0]        PE28_Out0;
wire [DWIDTH-1:0]        PE28_Out1;
wire [DWIDTH-1:0]        PE28_Out2;
wire [DWIDTH-1:0]        PE28_Out3;

wire [DWIDTH-1:0]        PE30_Out0;
wire [DWIDTH-1:0]        PE30_Out1;
wire [DWIDTH-1:0]        PE30_Out2;
wire [DWIDTH-1:0]        PE30_Out3;

wire [DWIDTH-1:0]        PE31_Out0;
wire [DWIDTH-1:0]        PE31_Out1;
wire [DWIDTH-1:0]        PE31_Out2;
wire [DWIDTH-1:0]        PE31_Out3;

wire [DWIDTH-1:0]        PE32_Out0;
wire [DWIDTH-1:0]        PE32_Out1;
wire [DWIDTH-1:0]        PE32_Out2;
wire [DWIDTH-1:0]        PE32_Out3;

wire [DWIDTH-1:0]        PE33_Out0;
wire [DWIDTH-1:0]        PE33_Out1;
wire [DWIDTH-1:0]        PE33_Out2;
wire [DWIDTH-1:0]        PE33_Out3;

wire [DWIDTH-1:0]        PE34_Out0;
wire [DWIDTH-1:0]        PE34_Out1;
wire [DWIDTH-1:0]        PE34_Out2;
wire [DWIDTH-1:0]        PE34_Out3;

wire [DWIDTH-1:0]        PE35_Out0;
wire [DWIDTH-1:0]        PE35_Out1;
wire [DWIDTH-1:0]        PE35_Out2;
wire [DWIDTH-1:0]        PE35_Out3;

wire [DWIDTH-1:0]        PE36_Out0;
wire [DWIDTH-1:0]        PE36_Out1;
wire [DWIDTH-1:0]        PE36_Out2;
wire [DWIDTH-1:0]        PE36_Out3;

wire [DWIDTH-1:0]        PE37_Out0;
wire [DWIDTH-1:0]        PE37_Out1;
wire [DWIDTH-1:0]        PE37_Out2;
wire [DWIDTH-1:0]        PE37_Out3;

wire [DWIDTH-1:0]        PE38_Out0;
wire [DWIDTH-1:0]        PE38_Out1;
wire [DWIDTH-1:0]        PE38_Out2;
wire [DWIDTH-1:0]        PE38_Out3;

wire [DWIDTH-1:0]        PE40_Out0;
wire [DWIDTH-1:0]        PE40_Out1;
wire [DWIDTH-1:0]        PE40_Out2;
wire [DWIDTH-1:0]        PE40_Out3;

wire [DWIDTH-1:0]        PE41_Out0;
wire [DWIDTH-1:0]        PE41_Out1;
wire [DWIDTH-1:0]        PE41_Out2;
wire [DWIDTH-1:0]        PE41_Out3;

wire [DWIDTH-1:0]        PE42_Out0;
wire [DWIDTH-1:0]        PE42_Out1;
wire [DWIDTH-1:0]        PE42_Out2;
wire [DWIDTH-1:0]        PE42_Out3;

wire [DWIDTH-1:0]        PE43_Out0;
wire [DWIDTH-1:0]        PE43_Out1;
wire [DWIDTH-1:0]        PE43_Out2;
wire [DWIDTH-1:0]        PE43_Out3;

wire [DWIDTH-1:0]        PE44_Out0;
wire [DWIDTH-1:0]        PE44_Out1;
wire [DWIDTH-1:0]        PE44_Out2;
wire [DWIDTH-1:0]        PE44_Out3;

wire [DWIDTH-1:0]        PE45_Out0;
wire [DWIDTH-1:0]        PE45_Out1;
wire [DWIDTH-1:0]        PE45_Out2;
wire [DWIDTH-1:0]        PE45_Out3;

wire [DWIDTH-1:0]        PE46_Out0;
wire [DWIDTH-1:0]        PE46_Out1;
wire [DWIDTH-1:0]        PE46_Out2;
wire [DWIDTH-1:0]        PE46_Out3;

wire [DWIDTH-1:0]        PE47_Out0;
wire [DWIDTH-1:0]        PE47_Out1;
wire [DWIDTH-1:0]        PE47_Out2;
wire [DWIDTH-1:0]        PE47_Out3;

wire [DWIDTH-1:0]        PE48_Out0;
wire [DWIDTH-1:0]        PE48_Out1;
wire [DWIDTH-1:0]        PE48_Out2;
wire [DWIDTH-1:0]        PE48_Out3;

wire [DWIDTH-1:0]        PE50_Out0;
wire [DWIDTH-1:0]        PE50_Out1;
wire [DWIDTH-1:0]        PE50_Out2;
wire [DWIDTH-1:0]        PE50_Out3;

wire [DWIDTH-1:0]        PE51_Out0;
wire [DWIDTH-1:0]        PE51_Out1;
wire [DWIDTH-1:0]        PE51_Out2;
wire [DWIDTH-1:0]        PE51_Out3;

wire [DWIDTH-1:0]        PE52_Out0;
wire [DWIDTH-1:0]        PE52_Out1;
wire [DWIDTH-1:0]        PE52_Out2;
wire [DWIDTH-1:0]        PE52_Out3;

wire [DWIDTH-1:0]        PE53_Out0;
wire [DWIDTH-1:0]        PE53_Out1;
wire [DWIDTH-1:0]        PE53_Out2;
wire [DWIDTH-1:0]        PE53_Out3;

wire [DWIDTH-1:0]        PE54_Out0;
wire [DWIDTH-1:0]        PE54_Out1;
wire [DWIDTH-1:0]        PE54_Out2;
wire [DWIDTH-1:0]        PE54_Out3;

wire [DWIDTH-1:0]        PE55_Out0;
wire [DWIDTH-1:0]        PE55_Out1;
wire [DWIDTH-1:0]        PE55_Out2;
wire [DWIDTH-1:0]        PE55_Out3;

wire [DWIDTH-1:0]        PE56_Out0;
wire [DWIDTH-1:0]        PE56_Out1;
wire [DWIDTH-1:0]        PE56_Out2;
wire [DWIDTH-1:0]        PE56_Out3;

wire [DWIDTH-1:0]        PE57_Out0;
wire [DWIDTH-1:0]        PE57_Out1;
wire [DWIDTH-1:0]        PE57_Out2;
wire [DWIDTH-1:0]        PE57_Out3;

wire [DWIDTH-1:0]        PE58_Out0;
wire [DWIDTH-1:0]        PE58_Out1;
wire [DWIDTH-1:0]        PE58_Out2;
wire [DWIDTH-1:0]        PE58_Out3;

wire [DWIDTH-1:0]        PE60_Out0;
wire [DWIDTH-1:0]        PE60_Out1;
wire [DWIDTH-1:0]        PE60_Out2;
wire [DWIDTH-1:0]        PE60_Out3;

wire [DWIDTH-1:0]        PE61_Out0;
wire [DWIDTH-1:0]        PE61_Out1;
wire [DWIDTH-1:0]        PE61_Out2;
wire [DWIDTH-1:0]        PE61_Out3;

wire [DWIDTH-1:0]        PE62_Out0;
wire [DWIDTH-1:0]        PE62_Out1;
wire [DWIDTH-1:0]        PE62_Out2;
wire [DWIDTH-1:0]        PE62_Out3;

wire [DWIDTH-1:0]        PE63_Out0;
wire [DWIDTH-1:0]        PE63_Out1;
wire [DWIDTH-1:0]        PE63_Out2;
wire [DWIDTH-1:0]        PE63_Out3;

wire [DWIDTH-1:0]        PE64_Out0;
wire [DWIDTH-1:0]        PE64_Out1;
wire [DWIDTH-1:0]        PE64_Out2;
wire [DWIDTH-1:0]        PE64_Out3;

wire [DWIDTH-1:0]        PE65_Out0;
wire [DWIDTH-1:0]        PE65_Out1;
wire [DWIDTH-1:0]        PE65_Out2;
wire [DWIDTH-1:0]        PE65_Out3;

wire [DWIDTH-1:0]        PE66_Out0;
wire [DWIDTH-1:0]        PE66_Out1;
wire [DWIDTH-1:0]        PE66_Out2;
wire [DWIDTH-1:0]        PE66_Out3;

wire [DWIDTH-1:0]        PE67_Out0;
wire [DWIDTH-1:0]        PE67_Out1;
wire [DWIDTH-1:0]        PE67_Out2;
wire [DWIDTH-1:0]        PE67_Out3;

wire [DWIDTH-1:0]        PE68_Out0;
wire [DWIDTH-1:0]        PE68_Out1;
wire [DWIDTH-1:0]        PE68_Out2;
wire [DWIDTH-1:0]        PE68_Out3;

wire [DWIDTH-1:0]        PE70_Out0;
wire [DWIDTH-1:0]        PE70_Out1;
wire [DWIDTH-1:0]        PE70_Out2;
wire [DWIDTH-1:0]        PE70_Out3;

wire [DWIDTH-1:0]        PE71_Out0;
wire [DWIDTH-1:0]        PE71_Out1;
wire [DWIDTH-1:0]        PE71_Out2;
wire [DWIDTH-1:0]        PE71_Out3;

wire [DWIDTH-1:0]        PE72_Out0;
wire [DWIDTH-1:0]        PE72_Out1;
wire [DWIDTH-1:0]        PE72_Out2;
wire [DWIDTH-1:0]        PE72_Out3;

wire [DWIDTH-1:0]        PE73_Out0;
wire [DWIDTH-1:0]        PE73_Out1;
wire [DWIDTH-1:0]        PE73_Out2;
wire [DWIDTH-1:0]        PE73_Out3;

wire [DWIDTH-1:0]        PE74_Out0;
wire [DWIDTH-1:0]        PE74_Out1;
wire [DWIDTH-1:0]        PE74_Out2;
wire [DWIDTH-1:0]        PE74_Out3;

wire [DWIDTH-1:0]        PE75_Out0;
wire [DWIDTH-1:0]        PE75_Out1;
wire [DWIDTH-1:0]        PE75_Out2;
wire [DWIDTH-1:0]        PE75_Out3;

wire [DWIDTH-1:0]        PE76_Out0;
wire [DWIDTH-1:0]        PE76_Out1;
wire [DWIDTH-1:0]        PE76_Out2;
wire [DWIDTH-1:0]        PE76_Out3;

wire [DWIDTH-1:0]        PE77_Out0;
wire [DWIDTH-1:0]        PE77_Out1;
wire [DWIDTH-1:0]        PE77_Out2;
wire [DWIDTH-1:0]        PE77_Out3;

wire [DWIDTH-1:0]        PE78_Out0;
wire [DWIDTH-1:0]        PE78_Out1;
wire [DWIDTH-1:0]        PE78_Out2;
wire [DWIDTH-1:0]        PE78_Out3;

wire [DWIDTH-1:0]        PE80_Out0;
wire [DWIDTH-1:0]        PE80_Out1;
wire [DWIDTH-1:0]        PE80_Out2;
wire [DWIDTH-1:0]        PE80_Out3;

wire [DWIDTH-1:0]        PE81_Out0;
wire [DWIDTH-1:0]        PE81_Out1;
wire [DWIDTH-1:0]        PE81_Out2;
wire [DWIDTH-1:0]        PE81_Out3;

wire [DWIDTH-1:0]        PE82_Out0;
wire [DWIDTH-1:0]        PE82_Out1;
wire [DWIDTH-1:0]        PE82_Out2;
wire [DWIDTH-1:0]        PE82_Out3;

wire [DWIDTH-1:0]        PE83_Out0;
wire [DWIDTH-1:0]        PE83_Out1;
wire [DWIDTH-1:0]        PE83_Out2;
wire [DWIDTH-1:0]        PE83_Out3;

wire [DWIDTH-1:0]        PE84_Out0;
wire [DWIDTH-1:0]        PE84_Out1;
wire [DWIDTH-1:0]        PE84_Out2;
wire [DWIDTH-1:0]        PE84_Out3;

wire [DWIDTH-1:0]        PE85_Out0;
wire [DWIDTH-1:0]        PE85_Out1;
wire [DWIDTH-1:0]        PE85_Out2;
wire [DWIDTH-1:0]        PE85_Out3;

wire [DWIDTH-1:0]        PE86_Out0;
wire [DWIDTH-1:0]        PE86_Out1;
wire [DWIDTH-1:0]        PE86_Out2;
wire [DWIDTH-1:0]        PE86_Out3;

wire [DWIDTH-1:0]        PE87_Out0;
wire [DWIDTH-1:0]        PE87_Out1;
wire [DWIDTH-1:0]        PE87_Out2;
wire [DWIDTH-1:0]        PE87_Out3;

wire [DWIDTH-1:0]        PE88_Out0;
wire [DWIDTH-1:0]        PE88_Out1;
wire [DWIDTH-1:0]        PE88_Out2;
wire [DWIDTH-1:0]        PE88_Out3;

wire [DWIDTH-1:0]        PE90_Out0;
wire [DWIDTH-1:0]        PE90_Out1;
wire [DWIDTH-1:0]        PE90_Out2;
wire [DWIDTH-1:0]        PE90_Out3;

wire [DWIDTH-1:0]        PE91_Out0;
wire [DWIDTH-1:0]        PE91_Out1;
wire [DWIDTH-1:0]        PE91_Out2;
wire [DWIDTH-1:0]        PE91_Out3;

wire [DWIDTH-1:0]        PE92_Out0;
wire [DWIDTH-1:0]        PE92_Out1;
wire [DWIDTH-1:0]        PE92_Out2;
wire [DWIDTH-1:0]        PE92_Out3;

wire [DWIDTH-1:0]        PE93_Out0;
wire [DWIDTH-1:0]        PE93_Out1;
wire [DWIDTH-1:0]        PE93_Out2;
wire [DWIDTH-1:0]        PE93_Out3;

wire [DWIDTH-1:0]        PE94_Out0;
wire [DWIDTH-1:0]        PE94_Out1;
wire [DWIDTH-1:0]        PE94_Out2;
wire [DWIDTH-1:0]        PE94_Out3;

wire [DWIDTH-1:0]        PE95_Out0;
wire [DWIDTH-1:0]        PE95_Out1;
wire [DWIDTH-1:0]        PE95_Out2;
wire [DWIDTH-1:0]        PE95_Out3;

wire [DWIDTH-1:0]        PE96_Out0;
wire [DWIDTH-1:0]        PE96_Out1;
wire [DWIDTH-1:0]        PE96_Out2;
wire [DWIDTH-1:0]        PE96_Out3;

wire [DWIDTH-1:0]        PE97_Out0;
wire [DWIDTH-1:0]        PE97_Out1;
wire [DWIDTH-1:0]        PE97_Out2;
wire [DWIDTH-1:0]        PE97_Out3;

wire [DWIDTH-1:0]        PE98_Out0;
wire [DWIDTH-1:0]        PE98_Out1;
wire [DWIDTH-1:0]        PE98_Out2;
wire [DWIDTH-1:0]        PE98_Out3;

PEIO PE00(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE08_Out2),
    .PE_In1(PE90_Out3),
    .PE_In2(PE01_Out0),
    .PE_In3(PE10_Out1),
    .PE_Out0(PE00_Out0),
    .PE_Out1(PE00_Out1),
    .PE_Out2(PE00_Out2),
    .PE_Out3(PE00_Out3),

    .PE_Load(Data0_Load),
    .PE_Store(Data0_Store),
    .PE_Array_Busy(PE_Array_Busy)

);
PEIO PE01(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE00_Out2),
    .PE_In1(PE91_Out3),
    .PE_In2(PE02_Out0),
    .PE_In3(PE11_Out1),
    .PE_Out0(PE01_Out0),
    .PE_Out1(PE01_Out1),
    .PE_Out2(PE01_Out2),
    .PE_Out3(PE01_Out3),

    .PE_Load(Data1_Load),
    .PE_Store(Data1_Store),
    .PE_Array_Busy(PE_Array_Busy)

);
PE PE02(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE01_Out2),
    .PE_In1(PE92_Out3),
    .PE_In2(PE03_Out0),
    .PE_In3(PE12_Out1),
    .PE_Out0(PE02_Out0),
    .PE_Out1(PE02_Out1),
    .PE_Out2(PE02_Out2),
    .PE_Out3(PE02_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE03(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE02_Out2),
    .PE_In1(PE93_Out3),
    .PE_In2(PE04_Out0),
    .PE_In3(PE13_Out1),
    .PE_Out0(PE03_Out0),
    .PE_Out1(PE03_Out1),
    .PE_Out2(PE03_Out2),
    .PE_Out3(PE03_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE04(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE03_Out2),
    .PE_In1(PE94_Out3),
    .PE_In2(PE05_Out0),
    .PE_In3(PE14_Out1),
    .PE_Out0(PE04_Out0),
    .PE_Out1(PE04_Out1),
    .PE_Out2(PE04_Out2),
    .PE_Out3(PE04_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE05(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE04_Out2),
    .PE_In1(PE95_Out3),
    .PE_In2(PE06_Out0),
    .PE_In3(PE15_Out1),
    .PE_Out0(PE05_Out0),
    .PE_Out1(PE05_Out1),
    .PE_Out2(PE05_Out2),
    .PE_Out3(PE05_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE06(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE05_Out2),
    .PE_In1(PE96_Out3),
    .PE_In2(PE07_Out0),
    .PE_In3(PE16_Out1),
    .PE_Out0(PE06_Out0),
    .PE_Out1(PE06_Out1),
    .PE_Out2(PE06_Out2),
    .PE_Out3(PE06_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE07(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE06_Out2),
    .PE_In1(PE97_Out3),
    .PE_In2(PE08_Out0),
    .PE_In3(PE17_Out1),
    .PE_Out0(PE07_Out0),
    .PE_Out1(PE07_Out1),
    .PE_Out2(PE07_Out2),
    .PE_Out3(PE07_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE08(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE07_Out2),
    .PE_In1(PE98_Out3),
    .PE_In2(PE00_Out0),
    .PE_In3(PE18_Out1),
    .PE_Out0(PE08_Out0),
    .PE_Out1(PE08_Out1),
    .PE_Out2(PE08_Out2),
    .PE_Out3(PE08_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE10(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE18_Out2),
    .PE_In1(PE00_Out3),
    .PE_In2(PE11_Out0),
    .PE_In3(PE20_Out1),
    .PE_Out0(PE10_Out0),
    .PE_Out1(PE10_Out1),
    .PE_Out2(PE10_Out2),
    .PE_Out3(PE10_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE11(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE10_Out2),
    .PE_In1(PE01_Out3),
    .PE_In2(PE12_Out0),
    .PE_In3(PE21_Out1),
    .PE_Out0(PE11_Out0),
    .PE_Out1(PE11_Out1),
    .PE_Out2(PE11_Out2),
    .PE_Out3(PE11_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE12(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE11_Out2),
    .PE_In1(PE02_Out3),
    .PE_In2(PE13_Out0),
    .PE_In3(PE22_Out1),
    .PE_Out0(PE12_Out0),
    .PE_Out1(PE12_Out1),
    .PE_Out2(PE12_Out2),
    .PE_Out3(PE12_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE13(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE12_Out2),
    .PE_In1(PE03_Out3),
    .PE_In2(PE14_Out0),
    .PE_In3(PE23_Out1),
    .PE_Out0(PE13_Out0),
    .PE_Out1(PE13_Out1),
    .PE_Out2(PE13_Out2),
    .PE_Out3(PE13_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE14(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE13_Out2),
    .PE_In1(PE04_Out3),
    .PE_In2(PE15_Out0),
    .PE_In3(PE24_Out1),
    .PE_Out0(PE14_Out0),
    .PE_Out1(PE14_Out1),
    .PE_Out2(PE14_Out2),
    .PE_Out3(PE14_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE15(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE14_Out2),
    .PE_In1(PE05_Out3),
    .PE_In2(PE16_Out0),
    .PE_In3(PE25_Out1),
    .PE_Out0(PE15_Out0),
    .PE_Out1(PE15_Out1),
    .PE_Out2(PE15_Out2),
    .PE_Out3(PE15_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE16(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE15_Out2),
    .PE_In1(PE06_Out3),
    .PE_In2(PE17_Out0),
    .PE_In3(PE26_Out1),
    .PE_Out0(PE16_Out0),
    .PE_Out1(PE16_Out1),
    .PE_Out2(PE16_Out2),
    .PE_Out3(PE16_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE17(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE16_Out2),
    .PE_In1(PE07_Out3),
    .PE_In2(PE18_Out0),
    .PE_In3(PE27_Out1),
    .PE_Out0(PE17_Out0),
    .PE_Out1(PE17_Out1),
    .PE_Out2(PE17_Out2),
    .PE_Out3(PE17_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE18(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE17_Out2),
    .PE_In1(PE08_Out3),
    .PE_In2(PE10_Out0),
    .PE_In3(PE28_Out1),
    .PE_Out0(PE18_Out0),
    .PE_Out1(PE18_Out1),
    .PE_Out2(PE18_Out2),
    .PE_Out3(PE18_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE20(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE28_Out2),
    .PE_In1(PE10_Out3),
    .PE_In2(PE21_Out0),
    .PE_In3(PE30_Out1),
    .PE_Out0(PE20_Out0),
    .PE_Out1(PE20_Out1),
    .PE_Out2(PE20_Out2),
    .PE_Out3(PE20_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE21(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE20_Out2),
    .PE_In1(PE11_Out3),
    .PE_In2(PE22_Out0),
    .PE_In3(PE31_Out1),
    .PE_Out0(PE21_Out0),
    .PE_Out1(PE21_Out1),
    .PE_Out2(PE21_Out2),
    .PE_Out3(PE21_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE22(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE21_Out2),
    .PE_In1(PE12_Out3),
    .PE_In2(PE23_Out0),
    .PE_In3(PE32_Out1),
    .PE_Out0(PE22_Out0),
    .PE_Out1(PE22_Out1),
    .PE_Out2(PE22_Out2),
    .PE_Out3(PE22_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE23(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE22_Out2),
    .PE_In1(PE13_Out3),
    .PE_In2(PE24_Out0),
    .PE_In3(PE33_Out1),
    .PE_Out0(PE23_Out0),
    .PE_Out1(PE23_Out1),
    .PE_Out2(PE23_Out2),
    .PE_Out3(PE23_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE24(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE23_Out2),
    .PE_In1(PE14_Out3),
    .PE_In2(PE25_Out0),
    .PE_In3(PE34_Out1),
    .PE_Out0(PE24_Out0),
    .PE_Out1(PE24_Out1),
    .PE_Out2(PE24_Out2),
    .PE_Out3(PE24_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE25(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE24_Out2),
    .PE_In1(PE15_Out3),
    .PE_In2(PE26_Out0),
    .PE_In3(PE35_Out1),
    .PE_Out0(PE25_Out0),
    .PE_Out1(PE25_Out1),
    .PE_Out2(PE25_Out2),
    .PE_Out3(PE25_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE26(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE25_Out2),
    .PE_In1(PE16_Out3),
    .PE_In2(PE27_Out0),
    .PE_In3(PE36_Out1),
    .PE_Out0(PE26_Out0),
    .PE_Out1(PE26_Out1),
    .PE_Out2(PE26_Out2),
    .PE_Out3(PE26_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE27(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE26_Out2),
    .PE_In1(PE17_Out3),
    .PE_In2(PE28_Out0),
    .PE_In3(PE37_Out1),
    .PE_Out0(PE27_Out0),
    .PE_Out1(PE27_Out1),
    .PE_Out2(PE27_Out2),
    .PE_Out3(PE27_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE28(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE27_Out2),
    .PE_In1(PE18_Out3),
    .PE_In2(PE20_Out0),
    .PE_In3(PE38_Out1),
    .PE_Out0(PE28_Out0),
    .PE_Out1(PE28_Out1),
    .PE_Out2(PE28_Out2),
    .PE_Out3(PE28_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE30(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE38_Out2),
    .PE_In1(PE20_Out3),
    .PE_In2(PE31_Out0),
    .PE_In3(PE40_Out1),
    .PE_Out0(PE30_Out0),
    .PE_Out1(PE30_Out1),
    .PE_Out2(PE30_Out2),
    .PE_Out3(PE30_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE31(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE30_Out2),
    .PE_In1(PE21_Out3),
    .PE_In2(PE32_Out0),
    .PE_In3(PE41_Out1),
    .PE_Out0(PE31_Out0),
    .PE_Out1(PE31_Out1),
    .PE_Out2(PE31_Out2),
    .PE_Out3(PE31_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE32(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE31_Out2),
    .PE_In1(PE22_Out3),
    .PE_In2(PE33_Out0),
    .PE_In3(PE42_Out1),
    .PE_Out0(PE32_Out0),
    .PE_Out1(PE32_Out1),
    .PE_Out2(PE32_Out2),
    .PE_Out3(PE32_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE33(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE32_Out2),
    .PE_In1(PE23_Out3),
    .PE_In2(PE34_Out0),
    .PE_In3(PE43_Out1),
    .PE_Out0(PE33_Out0),
    .PE_Out1(PE33_Out1),
    .PE_Out2(PE33_Out2),
    .PE_Out3(PE33_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE34(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE33_Out2),
    .PE_In1(PE24_Out3),
    .PE_In2(PE35_Out0),
    .PE_In3(PE44_Out1),
    .PE_Out0(PE34_Out0),
    .PE_Out1(PE34_Out1),
    .PE_Out2(PE34_Out2),
    .PE_Out3(PE34_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE35(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE34_Out2),
    .PE_In1(PE25_Out3),
    .PE_In2(PE36_Out0),
    .PE_In3(PE45_Out1),
    .PE_Out0(PE35_Out0),
    .PE_Out1(PE35_Out1),
    .PE_Out2(PE35_Out2),
    .PE_Out3(PE35_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE36(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE35_Out2),
    .PE_In1(PE26_Out3),
    .PE_In2(PE37_Out0),
    .PE_In3(PE46_Out1),
    .PE_Out0(PE36_Out0),
    .PE_Out1(PE36_Out1),
    .PE_Out2(PE36_Out2),
    .PE_Out3(PE36_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE37(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE36_Out2),
    .PE_In1(PE27_Out3),
    .PE_In2(PE38_Out0),
    .PE_In3(PE47_Out1),
    .PE_Out0(PE37_Out0),
    .PE_Out1(PE37_Out1),
    .PE_Out2(PE37_Out2),
    .PE_Out3(PE37_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE38(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE37_Out2),
    .PE_In1(PE28_Out3),
    .PE_In2(PE30_Out0),
    .PE_In3(PE48_Out1),
    .PE_Out0(PE38_Out0),
    .PE_Out1(PE38_Out1),
    .PE_Out2(PE38_Out2),
    .PE_Out3(PE38_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE40(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE48_Out2),
    .PE_In1(PE30_Out3),
    .PE_In2(PE41_Out0),
    .PE_In3(PE50_Out1),
    .PE_Out0(PE40_Out0),
    .PE_Out1(PE40_Out1),
    .PE_Out2(PE40_Out2),
    .PE_Out3(PE40_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE41(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE40_Out2),
    .PE_In1(PE31_Out3),
    .PE_In2(PE42_Out0),
    .PE_In3(PE51_Out1),
    .PE_Out0(PE41_Out0),
    .PE_Out1(PE41_Out1),
    .PE_Out2(PE41_Out2),
    .PE_Out3(PE41_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE42(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE41_Out2),
    .PE_In1(PE32_Out3),
    .PE_In2(PE43_Out0),
    .PE_In3(PE52_Out1),
    .PE_Out0(PE42_Out0),
    .PE_Out1(PE42_Out1),
    .PE_Out2(PE42_Out2),
    .PE_Out3(PE42_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE43(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE42_Out2),
    .PE_In1(PE33_Out3),
    .PE_In2(PE44_Out0),
    .PE_In3(PE53_Out1),
    .PE_Out0(PE43_Out0),
    .PE_Out1(PE43_Out1),
    .PE_Out2(PE43_Out2),
    .PE_Out3(PE43_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE44(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE43_Out2),
    .PE_In1(PE34_Out3),
    .PE_In2(PE45_Out0),
    .PE_In3(PE54_Out1),
    .PE_Out0(PE44_Out0),
    .PE_Out1(PE44_Out1),
    .PE_Out2(PE44_Out2),
    .PE_Out3(PE44_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE45(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE44_Out2),
    .PE_In1(PE35_Out3),
    .PE_In2(PE46_Out0),
    .PE_In3(PE55_Out1),
    .PE_Out0(PE45_Out0),
    .PE_Out1(PE45_Out1),
    .PE_Out2(PE45_Out2),
    .PE_Out3(PE45_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE46(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE45_Out2),
    .PE_In1(PE36_Out3),
    .PE_In2(PE47_Out0),
    .PE_In3(PE56_Out1),
    .PE_Out0(PE46_Out0),
    .PE_Out1(PE46_Out1),
    .PE_Out2(PE46_Out2),
    .PE_Out3(PE46_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE47(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE46_Out2),
    .PE_In1(PE37_Out3),
    .PE_In2(PE48_Out0),
    .PE_In3(PE57_Out1),
    .PE_Out0(PE47_Out0),
    .PE_Out1(PE47_Out1),
    .PE_Out2(PE47_Out2),
    .PE_Out3(PE47_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE48(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE47_Out2),
    .PE_In1(PE38_Out3),
    .PE_In2(PE40_Out0),
    .PE_In3(PE58_Out1),
    .PE_Out0(PE48_Out0),
    .PE_Out1(PE48_Out1),
    .PE_Out2(PE48_Out2),
    .PE_Out3(PE48_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE50(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE58_Out2),
    .PE_In1(PE40_Out3),
    .PE_In2(PE51_Out0),
    .PE_In3(PE60_Out1),
    .PE_Out0(PE50_Out0),
    .PE_Out1(PE50_Out1),
    .PE_Out2(PE50_Out2),
    .PE_Out3(PE50_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE51(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE50_Out2),
    .PE_In1(PE41_Out3),
    .PE_In2(PE52_Out0),
    .PE_In3(PE61_Out1),
    .PE_Out0(PE51_Out0),
    .PE_Out1(PE51_Out1),
    .PE_Out2(PE51_Out2),
    .PE_Out3(PE51_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE52(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE51_Out2),
    .PE_In1(PE42_Out3),
    .PE_In2(PE53_Out0),
    .PE_In3(PE62_Out1),
    .PE_Out0(PE52_Out0),
    .PE_Out1(PE52_Out1),
    .PE_Out2(PE52_Out2),
    .PE_Out3(PE52_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE53(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE52_Out2),
    .PE_In1(PE43_Out3),
    .PE_In2(PE54_Out0),
    .PE_In3(PE63_Out1),
    .PE_Out0(PE53_Out0),
    .PE_Out1(PE53_Out1),
    .PE_Out2(PE53_Out2),
    .PE_Out3(PE53_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE54(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE53_Out2),
    .PE_In1(PE44_Out3),
    .PE_In2(PE55_Out0),
    .PE_In3(PE64_Out1),
    .PE_Out0(PE54_Out0),
    .PE_Out1(PE54_Out1),
    .PE_Out2(PE54_Out2),
    .PE_Out3(PE54_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE55(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE54_Out2),
    .PE_In1(PE45_Out3),
    .PE_In2(PE56_Out0),
    .PE_In3(PE65_Out1),
    .PE_Out0(PE55_Out0),
    .PE_Out1(PE55_Out1),
    .PE_Out2(PE55_Out2),
    .PE_Out3(PE55_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE56(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE55_Out2),
    .PE_In1(PE46_Out3),
    .PE_In2(PE57_Out0),
    .PE_In3(PE66_Out1),
    .PE_Out0(PE56_Out0),
    .PE_Out1(PE56_Out1),
    .PE_Out2(PE56_Out2),
    .PE_Out3(PE56_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE57(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE56_Out2),
    .PE_In1(PE47_Out3),
    .PE_In2(PE58_Out0),
    .PE_In3(PE67_Out1),
    .PE_Out0(PE57_Out0),
    .PE_Out1(PE57_Out1),
    .PE_Out2(PE57_Out2),
    .PE_Out3(PE57_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE58(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE57_Out2),
    .PE_In1(PE48_Out3),
    .PE_In2(PE50_Out0),
    .PE_In3(PE68_Out1),
    .PE_Out0(PE58_Out0),
    .PE_Out1(PE58_Out1),
    .PE_Out2(PE58_Out2),
    .PE_Out3(PE58_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE60(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE68_Out2),
    .PE_In1(PE50_Out3),
    .PE_In2(PE61_Out0),
    .PE_In3(PE70_Out1),
    .PE_Out0(PE60_Out0),
    .PE_Out1(PE60_Out1),
    .PE_Out2(PE60_Out2),
    .PE_Out3(PE60_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE61(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE60_Out2),
    .PE_In1(PE51_Out3),
    .PE_In2(PE62_Out0),
    .PE_In3(PE71_Out1),
    .PE_Out0(PE61_Out0),
    .PE_Out1(PE61_Out1),
    .PE_Out2(PE61_Out2),
    .PE_Out3(PE61_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE62(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE61_Out2),
    .PE_In1(PE52_Out3),
    .PE_In2(PE63_Out0),
    .PE_In3(PE72_Out1),
    .PE_Out0(PE62_Out0),
    .PE_Out1(PE62_Out1),
    .PE_Out2(PE62_Out2),
    .PE_Out3(PE62_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE63(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE62_Out2),
    .PE_In1(PE53_Out3),
    .PE_In2(PE64_Out0),
    .PE_In3(PE73_Out1),
    .PE_Out0(PE63_Out0),
    .PE_Out1(PE63_Out1),
    .PE_Out2(PE63_Out2),
    .PE_Out3(PE63_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE64(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE63_Out2),
    .PE_In1(PE54_Out3),
    .PE_In2(PE65_Out0),
    .PE_In3(PE74_Out1),
    .PE_Out0(PE64_Out0),
    .PE_Out1(PE64_Out1),
    .PE_Out2(PE64_Out2),
    .PE_Out3(PE64_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE65(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE64_Out2),
    .PE_In1(PE55_Out3),
    .PE_In2(PE66_Out0),
    .PE_In3(PE75_Out1),
    .PE_Out0(PE65_Out0),
    .PE_Out1(PE65_Out1),
    .PE_Out2(PE65_Out2),
    .PE_Out3(PE65_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE66(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE65_Out2),
    .PE_In1(PE56_Out3),
    .PE_In2(PE67_Out0),
    .PE_In3(PE76_Out1),
    .PE_Out0(PE66_Out0),
    .PE_Out1(PE66_Out1),
    .PE_Out2(PE66_Out2),
    .PE_Out3(PE66_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE67(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE66_Out2),
    .PE_In1(PE57_Out3),
    .PE_In2(PE68_Out0),
    .PE_In3(PE77_Out1),
    .PE_Out0(PE67_Out0),
    .PE_Out1(PE67_Out1),
    .PE_Out2(PE67_Out2),
    .PE_Out3(PE67_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE68(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE67_Out2),
    .PE_In1(PE58_Out3),
    .PE_In2(PE60_Out0),
    .PE_In3(PE78_Out1),
    .PE_Out0(PE68_Out0),
    .PE_Out1(PE68_Out1),
    .PE_Out2(PE68_Out2),
    .PE_Out3(PE68_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE70(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE78_Out2),
    .PE_In1(PE60_Out3),
    .PE_In2(PE71_Out0),
    .PE_In3(PE80_Out1),
    .PE_Out0(PE70_Out0),
    .PE_Out1(PE70_Out1),
    .PE_Out2(PE70_Out2),
    .PE_Out3(PE70_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE71(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE70_Out2),
    .PE_In1(PE61_Out3),
    .PE_In2(PE72_Out0),
    .PE_In3(PE81_Out1),
    .PE_Out0(PE71_Out0),
    .PE_Out1(PE71_Out1),
    .PE_Out2(PE71_Out2),
    .PE_Out3(PE71_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE72(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE71_Out2),
    .PE_In1(PE62_Out3),
    .PE_In2(PE73_Out0),
    .PE_In3(PE82_Out1),
    .PE_Out0(PE72_Out0),
    .PE_Out1(PE72_Out1),
    .PE_Out2(PE72_Out2),
    .PE_Out3(PE72_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE73(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE72_Out2),
    .PE_In1(PE63_Out3),
    .PE_In2(PE74_Out0),
    .PE_In3(PE83_Out1),
    .PE_Out0(PE73_Out0),
    .PE_Out1(PE73_Out1),
    .PE_Out2(PE73_Out2),
    .PE_Out3(PE73_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE74(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE73_Out2),
    .PE_In1(PE64_Out3),
    .PE_In2(PE75_Out0),
    .PE_In3(PE84_Out1),
    .PE_Out0(PE74_Out0),
    .PE_Out1(PE74_Out1),
    .PE_Out2(PE74_Out2),
    .PE_Out3(PE74_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE75(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE74_Out2),
    .PE_In1(PE65_Out3),
    .PE_In2(PE76_Out0),
    .PE_In3(PE85_Out1),
    .PE_Out0(PE75_Out0),
    .PE_Out1(PE75_Out1),
    .PE_Out2(PE75_Out2),
    .PE_Out3(PE75_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE76(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE75_Out2),
    .PE_In1(PE66_Out3),
    .PE_In2(PE77_Out0),
    .PE_In3(PE86_Out1),
    .PE_Out0(PE76_Out0),
    .PE_Out1(PE76_Out1),
    .PE_Out2(PE76_Out2),
    .PE_Out3(PE76_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE77(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE76_Out2),
    .PE_In1(PE67_Out3),
    .PE_In2(PE78_Out0),
    .PE_In3(PE87_Out1),
    .PE_Out0(PE77_Out0),
    .PE_Out1(PE77_Out1),
    .PE_Out2(PE77_Out2),
    .PE_Out3(PE77_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE78(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE77_Out2),
    .PE_In1(PE68_Out3),
    .PE_In2(PE70_Out0),
    .PE_In3(PE88_Out1),
    .PE_Out0(PE78_Out0),
    .PE_Out1(PE78_Out1),
    .PE_Out2(PE78_Out2),
    .PE_Out3(PE78_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE80(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE88_Out2),
    .PE_In1(PE70_Out3),
    .PE_In2(PE81_Out0),
    .PE_In3(PE90_Out1),
    .PE_Out0(PE80_Out0),
    .PE_Out1(PE80_Out1),
    .PE_Out2(PE80_Out2),
    .PE_Out3(PE80_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE81(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE80_Out2),
    .PE_In1(PE71_Out3),
    .PE_In2(PE82_Out0),
    .PE_In3(PE91_Out1),
    .PE_Out0(PE81_Out0),
    .PE_Out1(PE81_Out1),
    .PE_Out2(PE81_Out2),
    .PE_Out3(PE81_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE82(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE81_Out2),
    .PE_In1(PE72_Out3),
    .PE_In2(PE83_Out0),
    .PE_In3(PE92_Out1),
    .PE_Out0(PE82_Out0),
    .PE_Out1(PE82_Out1),
    .PE_Out2(PE82_Out2),
    .PE_Out3(PE82_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE83(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE82_Out2),
    .PE_In1(PE73_Out3),
    .PE_In2(PE84_Out0),
    .PE_In3(PE93_Out1),
    .PE_Out0(PE83_Out0),
    .PE_Out1(PE83_Out1),
    .PE_Out2(PE83_Out2),
    .PE_Out3(PE83_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE84(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE83_Out2),
    .PE_In1(PE74_Out3),
    .PE_In2(PE85_Out0),
    .PE_In3(PE94_Out1),
    .PE_Out0(PE84_Out0),
    .PE_Out1(PE84_Out1),
    .PE_Out2(PE84_Out2),
    .PE_Out3(PE84_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE85(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE84_Out2),
    .PE_In1(PE75_Out3),
    .PE_In2(PE86_Out0),
    .PE_In3(PE95_Out1),
    .PE_Out0(PE85_Out0),
    .PE_Out1(PE85_Out1),
    .PE_Out2(PE85_Out2),
    .PE_Out3(PE85_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE86(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE85_Out2),
    .PE_In1(PE76_Out3),
    .PE_In2(PE87_Out0),
    .PE_In3(PE96_Out1),
    .PE_Out0(PE86_Out0),
    .PE_Out1(PE86_Out1),
    .PE_Out2(PE86_Out2),
    .PE_Out3(PE86_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE87(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE86_Out2),
    .PE_In1(PE77_Out3),
    .PE_In2(PE88_Out0),
    .PE_In3(PE97_Out1),
    .PE_Out0(PE87_Out0),
    .PE_Out1(PE87_Out1),
    .PE_Out2(PE87_Out2),
    .PE_Out3(PE87_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE88(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE87_Out2),
    .PE_In1(PE78_Out3),
    .PE_In2(PE80_Out0),
    .PE_In3(PE98_Out1),
    .PE_Out0(PE88_Out0),
    .PE_Out1(PE88_Out1),
    .PE_Out2(PE88_Out2),
    .PE_Out3(PE88_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE90(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE98_Out2),
    .PE_In1(PE80_Out3),
    .PE_In2(PE91_Out0),
    .PE_In3(PE00_Out1),
    .PE_Out0(PE90_Out0),
    .PE_Out1(PE90_Out1),
    .PE_Out2(PE90_Out2),
    .PE_Out3(PE90_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE91(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE90_Out2),
    .PE_In1(PE81_Out3),
    .PE_In2(PE92_Out0),
    .PE_In3(PE01_Out1),
    .PE_Out0(PE91_Out0),
    .PE_Out1(PE91_Out1),
    .PE_Out2(PE91_Out2),
    .PE_Out3(PE91_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE92(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE91_Out2),
    .PE_In1(PE82_Out3),
    .PE_In2(PE93_Out0),
    .PE_In3(PE02_Out1),
    .PE_Out0(PE92_Out0),
    .PE_Out1(PE92_Out1),
    .PE_Out2(PE92_Out2),
    .PE_Out3(PE92_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE93(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE92_Out2),
    .PE_In1(PE83_Out3),
    .PE_In2(PE94_Out0),
    .PE_In3(PE03_Out1),
    .PE_Out0(PE93_Out0),
    .PE_Out1(PE93_Out1),
    .PE_Out2(PE93_Out2),
    .PE_Out3(PE93_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE94(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE93_Out2),
    .PE_In1(PE84_Out3),
    .PE_In2(PE95_Out0),
    .PE_In3(PE04_Out1),
    .PE_Out0(PE94_Out0),
    .PE_Out1(PE94_Out1),
    .PE_Out2(PE94_Out2),
    .PE_Out3(PE94_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE95(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE94_Out2),
    .PE_In1(PE85_Out3),
    .PE_In2(PE96_Out0),
    .PE_In3(PE05_Out1),
    .PE_Out0(PE95_Out0),
    .PE_Out1(PE95_Out1),
    .PE_Out2(PE95_Out2),
    .PE_Out3(PE95_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE96(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE95_Out2),
    .PE_In1(PE86_Out3),
    .PE_In2(PE97_Out0),
    .PE_In3(PE06_Out1),
    .PE_Out0(PE96_Out0),
    .PE_Out1(PE96_Out1),
    .PE_Out2(PE96_Out2),
    .PE_Out3(PE96_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE97(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE96_Out2),
    .PE_In1(PE87_Out3),
    .PE_In2(PE98_Out0),
    .PE_In3(PE07_Out1),
    .PE_Out0(PE97_Out0),
    .PE_Out1(PE97_Out1),
    .PE_Out2(PE97_Out2),
    .PE_Out3(PE97_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE98(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE97_Out2),
    .PE_In1(PE88_Out3),
    .PE_In2(PE90_Out0),
    .PE_In3(PE08_Out1),
    .PE_Out0(PE98_Out0),
    .PE_Out1(PE98_Out1),
    .PE_Out2(PE98_Out2),
    .PE_Out3(PE98_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
endmodule
