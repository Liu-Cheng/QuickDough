`timescale 1ns / 1ps

module torus128(
	      clk,
          rst_n,
          data_out0,
          data_out1,
          data_out2,
          data_out3
	      );

input clk;
input rst_n;

output[15:0] data_out0;
output[15:0] data_out1;
output[15:0] data_out2;
output[15:0] data_out3;

wire [15:0] PE00_out0;
wire [15:0] PE00_out1;
wire [15:0] PE00_out2;
wire [15:0] PE00_out3;

wire [15:0] PE01_out0;
wire [15:0] PE01_out1;
wire [15:0] PE01_out2;
wire [15:0] PE01_out3;

wire [15:0] PE02_out0;
wire [15:0] PE02_out1;
wire [15:0] PE02_out2;
wire [15:0] PE02_out3;

wire [15:0] PE03_out0;
wire [15:0] PE03_out1;
wire [15:0] PE03_out2;
wire [15:0] PE03_out3;

wire [15:0] PE04_out0;
wire [15:0] PE04_out1;
wire [15:0] PE04_out2;
wire [15:0] PE04_out3;

wire [15:0] PE05_out0;
wire [15:0] PE05_out1;
wire [15:0] PE05_out2;
wire [15:0] PE05_out3;

wire [15:0] PE06_out0;
wire [15:0] PE06_out1;
wire [15:0] PE06_out2;
wire [15:0] PE06_out3;

wire [15:0] PE07_out0;
wire [15:0] PE07_out1;
wire [15:0] PE07_out2;
wire [15:0] PE07_out3;


wire [15:0] PE10_out0;
wire [15:0] PE10_out1;
wire [15:0] PE10_out2;
wire [15:0] PE10_out3;

wire [15:0] PE11_out0;
wire [15:0] PE11_out1;
wire [15:0] PE11_out2;
wire [15:0] PE11_out3;

wire [15:0] PE12_out0;
wire [15:0] PE12_out1;
wire [15:0] PE12_out2;
wire [15:0] PE12_out3;

wire [15:0] PE13_out0;
wire [15:0] PE13_out1;
wire [15:0] PE13_out2;
wire [15:0] PE13_out3;

wire [15:0] PE14_out0;
wire [15:0] PE14_out1;
wire [15:0] PE14_out2;
wire [15:0] PE14_out3;

wire [15:0] PE15_out0;
wire [15:0] PE15_out1;
wire [15:0] PE15_out2;
wire [15:0] PE15_out3;

wire [15:0] PE16_out0;
wire [15:0] PE16_out1;
wire [15:0] PE16_out2;
wire [15:0] PE16_out3;

wire [15:0] PE17_out0;
wire [15:0] PE17_out1;
wire [15:0] PE17_out2;
wire [15:0] PE17_out3;


wire [15:0] PE20_out0;
wire [15:0] PE20_out1;
wire [15:0] PE20_out2;
wire [15:0] PE20_out3;

wire [15:0] PE21_out0;
wire [15:0] PE21_out1;
wire [15:0] PE21_out2;
wire [15:0] PE21_out3;

wire [15:0] PE22_out0;
wire [15:0] PE22_out1;
wire [15:0] PE22_out2;
wire [15:0] PE22_out3;

wire [15:0] PE23_out0;
wire [15:0] PE23_out1;
wire [15:0] PE23_out2;
wire [15:0] PE23_out3;

wire [15:0] PE24_out0;
wire [15:0] PE24_out1;
wire [15:0] PE24_out2;
wire [15:0] PE24_out3;

wire [15:0] PE25_out0;
wire [15:0] PE25_out1;
wire [15:0] PE25_out2;
wire [15:0] PE25_out3;

wire [15:0] PE26_out0;
wire [15:0] PE26_out1;
wire [15:0] PE26_out2;
wire [15:0] PE26_out3;

wire [15:0] PE27_out0;
wire [15:0] PE27_out1;
wire [15:0] PE27_out2;
wire [15:0] PE27_out3;


wire [15:0] PE30_out0;
wire [15:0] PE30_out1;
wire [15:0] PE30_out2;
wire [15:0] PE30_out3;

wire [15:0] PE31_out0;
wire [15:0] PE31_out1;
wire [15:0] PE31_out2;
wire [15:0] PE31_out3;

wire [15:0] PE32_out0;
wire [15:0] PE32_out1;
wire [15:0] PE32_out2;
wire [15:0] PE32_out3;

wire [15:0] PE33_out0;
wire [15:0] PE33_out1;
wire [15:0] PE33_out2;
wire [15:0] PE33_out3;

wire [15:0] PE34_out0;
wire [15:0] PE34_out1;
wire [15:0] PE34_out2;
wire [15:0] PE34_out3;

wire [15:0] PE35_out0;
wire [15:0] PE35_out1;
wire [15:0] PE35_out2;
wire [15:0] PE35_out3;

wire [15:0] PE36_out0;
wire [15:0] PE36_out1;
wire [15:0] PE36_out2;
wire [15:0] PE36_out3;

wire [15:0] PE37_out0;
wire [15:0] PE37_out1;
wire [15:0] PE37_out2;
wire [15:0] PE37_out3;


wire [15:0] PE40_out0;
wire [15:0] PE40_out1;
wire [15:0] PE40_out2;
wire [15:0] PE40_out3;

wire [15:0] PE41_out0;
wire [15:0] PE41_out1;
wire [15:0] PE41_out2;
wire [15:0] PE41_out3;

wire [15:0] PE42_out0;
wire [15:0] PE42_out1;
wire [15:0] PE42_out2;
wire [15:0] PE42_out3;

wire [15:0] PE43_out0;
wire [15:0] PE43_out1;
wire [15:0] PE43_out2;
wire [15:0] PE43_out3;

wire [15:0] PE44_out0;
wire [15:0] PE44_out1;
wire [15:0] PE44_out2;
wire [15:0] PE44_out3;

wire [15:0] PE45_out0;
wire [15:0] PE45_out1;
wire [15:0] PE45_out2;
wire [15:0] PE45_out3;

wire [15:0] PE46_out0;
wire [15:0] PE46_out1;
wire [15:0] PE46_out2;
wire [15:0] PE46_out3;

wire [15:0] PE47_out0;
wire [15:0] PE47_out1;
wire [15:0] PE47_out2;
wire [15:0] PE47_out3;


wire [15:0] PE50_out0;
wire [15:0] PE50_out1;
wire [15:0] PE50_out2;
wire [15:0] PE50_out3;

wire [15:0] PE51_out0;
wire [15:0] PE51_out1;
wire [15:0] PE51_out2;
wire [15:0] PE51_out3;

wire [15:0] PE52_out0;
wire [15:0] PE52_out1;
wire [15:0] PE52_out2;
wire [15:0] PE52_out3;

wire [15:0] PE53_out0;
wire [15:0] PE53_out1;
wire [15:0] PE53_out2;
wire [15:0] PE53_out3;

wire [15:0] PE54_out0;
wire [15:0] PE54_out1;
wire [15:0] PE54_out2;
wire [15:0] PE54_out3;

wire [15:0] PE55_out0;
wire [15:0] PE55_out1;
wire [15:0] PE55_out2;
wire [15:0] PE55_out3;

wire [15:0] PE56_out0;
wire [15:0] PE56_out1;
wire [15:0] PE56_out2;
wire [15:0] PE56_out3;

wire [15:0] PE57_out0;
wire [15:0] PE57_out1;
wire [15:0] PE57_out2;
wire [15:0] PE57_out3;


wire [15:0] PE60_out0;
wire [15:0] PE60_out1;
wire [15:0] PE60_out2;
wire [15:0] PE60_out3;

wire [15:0] PE61_out0;
wire [15:0] PE61_out1;
wire [15:0] PE61_out2;
wire [15:0] PE61_out3;

wire [15:0] PE62_out0;
wire [15:0] PE62_out1;
wire [15:0] PE62_out2;
wire [15:0] PE62_out3;

wire [15:0] PE63_out0;
wire [15:0] PE63_out1;
wire [15:0] PE63_out2;
wire [15:0] PE63_out3;

wire [15:0] PE64_out0;
wire [15:0] PE64_out1;
wire [15:0] PE64_out2;
wire [15:0] PE64_out3;

wire [15:0] PE65_out0;
wire [15:0] PE65_out1;
wire [15:0] PE65_out2;
wire [15:0] PE65_out3;

wire [15:0] PE66_out0;
wire [15:0] PE66_out1;
wire [15:0] PE66_out2;
wire [15:0] PE66_out3;

wire [15:0] PE67_out0;
wire [15:0] PE67_out1;
wire [15:0] PE67_out2;
wire [15:0] PE67_out3;


wire [15:0] PE70_out0;
wire [15:0] PE70_out1;
wire [15:0] PE70_out2;
wire [15:0] PE70_out3;

wire [15:0] PE71_out0;
wire [15:0] PE71_out1;
wire [15:0] PE71_out2;
wire [15:0] PE71_out3;

wire [15:0] PE72_out0;
wire [15:0] PE72_out1;
wire [15:0] PE72_out2;
wire [15:0] PE72_out3;

wire [15:0] PE73_out0;
wire [15:0] PE73_out1;
wire [15:0] PE73_out2;
wire [15:0] PE73_out3;

wire [15:0] PE74_out0;
wire [15:0] PE74_out1;
wire [15:0] PE74_out2;
wire [15:0] PE74_out3;

wire [15:0] PE75_out0;
wire [15:0] PE75_out1;
wire [15:0] PE75_out2;
wire [15:0] PE75_out3;

wire [15:0] PE76_out0;
wire [15:0] PE76_out1;
wire [15:0] PE76_out2;
wire [15:0] PE76_out3;

wire [15:0] PE77_out0;
wire [15:0] PE77_out1;
wire [15:0] PE77_out2;
wire [15:0] PE77_out3;


wire [15:0] PE80_out0;
wire [15:0] PE80_out1;
wire [15:0] PE80_out2;
wire [15:0] PE80_out3;

wire [15:0] PE81_out0;
wire [15:0] PE81_out1;
wire [15:0] PE81_out2;
wire [15:0] PE81_out3;

wire [15:0] PE82_out0;
wire [15:0] PE82_out1;
wire [15:0] PE82_out2;
wire [15:0] PE82_out3;

wire [15:0] PE83_out0;
wire [15:0] PE83_out1;
wire [15:0] PE83_out2;
wire [15:0] PE83_out3;

wire [15:0] PE84_out0;
wire [15:0] PE84_out1;
wire [15:0] PE84_out2;
wire [15:0] PE84_out3;

wire [15:0] PE85_out0;
wire [15:0] PE85_out1;
wire [15:0] PE85_out2;
wire [15:0] PE85_out3;

wire [15:0] PE86_out0;
wire [15:0] PE86_out1;
wire [15:0] PE86_out2;
wire [15:0] PE86_out3;

wire [15:0] PE87_out0;
wire [15:0] PE87_out1;
wire [15:0] PE87_out2;
wire [15:0] PE87_out3;


wire [15:0] PE90_out0;
wire [15:0] PE90_out1;
wire [15:0] PE90_out2;
wire [15:0] PE90_out3;

wire [15:0] PE91_out0;
wire [15:0] PE91_out1;
wire [15:0] PE91_out2;
wire [15:0] PE91_out3;

wire [15:0] PE92_out0;
wire [15:0] PE92_out1;
wire [15:0] PE92_out2;
wire [15:0] PE92_out3;

wire [15:0] PE93_out0;
wire [15:0] PE93_out1;
wire [15:0] PE93_out2;
wire [15:0] PE93_out3;

wire [15:0] PE94_out0;
wire [15:0] PE94_out1;
wire [15:0] PE94_out2;
wire [15:0] PE94_out3;

wire [15:0] PE95_out0;
wire [15:0] PE95_out1;
wire [15:0] PE95_out2;
wire [15:0] PE95_out3;

wire [15:0] PE96_out0;
wire [15:0] PE96_out1;
wire [15:0] PE96_out2;
wire [15:0] PE96_out3;

wire [15:0] PE97_out0;
wire [15:0] PE97_out1;
wire [15:0] PE97_out2;
wire [15:0] PE97_out3;


wire [15:0] PE100_out0;
wire [15:0] PE100_out1;
wire [15:0] PE100_out2;
wire [15:0] PE100_out3;

wire [15:0] PE101_out0;
wire [15:0] PE101_out1;
wire [15:0] PE101_out2;
wire [15:0] PE101_out3;

wire [15:0] PE102_out0;
wire [15:0] PE102_out1;
wire [15:0] PE102_out2;
wire [15:0] PE102_out3;

wire [15:0] PE103_out0;
wire [15:0] PE103_out1;
wire [15:0] PE103_out2;
wire [15:0] PE103_out3;

wire [15:0] PE104_out0;
wire [15:0] PE104_out1;
wire [15:0] PE104_out2;
wire [15:0] PE104_out3;

wire [15:0] PE105_out0;
wire [15:0] PE105_out1;
wire [15:0] PE105_out2;
wire [15:0] PE105_out3;

wire [15:0] PE106_out0;
wire [15:0] PE106_out1;
wire [15:0] PE106_out2;
wire [15:0] PE106_out3;

wire [15:0] PE107_out0;
wire [15:0] PE107_out1;
wire [15:0] PE107_out2;
wire [15:0] PE107_out3;


wire [15:0] PE110_out0;
wire [15:0] PE110_out1;
wire [15:0] PE110_out2;
wire [15:0] PE110_out3;

wire [15:0] PE111_out0;
wire [15:0] PE111_out1;
wire [15:0] PE111_out2;
wire [15:0] PE111_out3;

wire [15:0] PE112_out0;
wire [15:0] PE112_out1;
wire [15:0] PE112_out2;
wire [15:0] PE112_out3;

wire [15:0] PE113_out0;
wire [15:0] PE113_out1;
wire [15:0] PE113_out2;
wire [15:0] PE113_out3;

wire [15:0] PE114_out0;
wire [15:0] PE114_out1;
wire [15:0] PE114_out2;
wire [15:0] PE114_out3;

wire [15:0] PE115_out0;
wire [15:0] PE115_out1;
wire [15:0] PE115_out2;
wire [15:0] PE115_out3;

wire [15:0] PE116_out0;
wire [15:0] PE116_out1;
wire [15:0] PE116_out2;
wire [15:0] PE116_out3;

wire [15:0] PE117_out0;
wire [15:0] PE117_out1;
wire [15:0] PE117_out2;
wire [15:0] PE117_out3;


wire [15:0] PE120_out0;
wire [15:0] PE120_out1;
wire [15:0] PE120_out2;
wire [15:0] PE120_out3;

wire [15:0] PE121_out0;
wire [15:0] PE121_out1;
wire [15:0] PE121_out2;
wire [15:0] PE121_out3;

wire [15:0] PE122_out0;
wire [15:0] PE122_out1;
wire [15:0] PE122_out2;
wire [15:0] PE122_out3;

wire [15:0] PE123_out0;
wire [15:0] PE123_out1;
wire [15:0] PE123_out2;
wire [15:0] PE123_out3;

wire [15:0] PE124_out0;
wire [15:0] PE124_out1;
wire [15:0] PE124_out2;
wire [15:0] PE124_out3;

wire [15:0] PE125_out0;
wire [15:0] PE125_out1;
wire [15:0] PE125_out2;
wire [15:0] PE125_out3;

wire [15:0] PE126_out0;
wire [15:0] PE126_out1;
wire [15:0] PE126_out2;
wire [15:0] PE126_out3;

wire [15:0] PE127_out0;
wire [15:0] PE127_out1;
wire [15:0] PE127_out2;
wire [15:0] PE127_out3;


wire [15:0] PE130_out0;
wire [15:0] PE130_out1;
wire [15:0] PE130_out2;
wire [15:0] PE130_out3;

wire [15:0] PE131_out0;
wire [15:0] PE131_out1;
wire [15:0] PE131_out2;
wire [15:0] PE131_out3;

wire [15:0] PE132_out0;
wire [15:0] PE132_out1;
wire [15:0] PE132_out2;
wire [15:0] PE132_out3;

wire [15:0] PE133_out0;
wire [15:0] PE133_out1;
wire [15:0] PE133_out2;
wire [15:0] PE133_out3;

wire [15:0] PE134_out0;
wire [15:0] PE134_out1;
wire [15:0] PE134_out2;
wire [15:0] PE134_out3;

wire [15:0] PE135_out0;
wire [15:0] PE135_out1;
wire [15:0] PE135_out2;
wire [15:0] PE135_out3;

wire [15:0] PE136_out0;
wire [15:0] PE136_out1;
wire [15:0] PE136_out2;
wire [15:0] PE136_out3;

wire [15:0] PE137_out0;
wire [15:0] PE137_out1;
wire [15:0] PE137_out2;
wire [15:0] PE137_out3;


wire [15:0] PE140_out0;
wire [15:0] PE140_out1;
wire [15:0] PE140_out2;
wire [15:0] PE140_out3;

wire [15:0] PE141_out0;
wire [15:0] PE141_out1;
wire [15:0] PE141_out2;
wire [15:0] PE141_out3;

wire [15:0] PE142_out0;
wire [15:0] PE142_out1;
wire [15:0] PE142_out2;
wire [15:0] PE142_out3;

wire [15:0] PE143_out0;
wire [15:0] PE143_out1;
wire [15:0] PE143_out2;
wire [15:0] PE143_out3;

wire [15:0] PE144_out0;
wire [15:0] PE144_out1;
wire [15:0] PE144_out2;
wire [15:0] PE144_out3;

wire [15:0] PE145_out0;
wire [15:0] PE145_out1;
wire [15:0] PE145_out2;
wire [15:0] PE145_out3;

wire [15:0] PE146_out0;
wire [15:0] PE146_out1;
wire [15:0] PE146_out2;
wire [15:0] PE146_out3;

wire [15:0] PE147_out0;
wire [15:0] PE147_out1;
wire [15:0] PE147_out2;
wire [15:0] PE147_out3;


wire [15:0] PE150_out0;
wire [15:0] PE150_out1;
wire [15:0] PE150_out2;
wire [15:0] PE150_out3;

wire [15:0] PE151_out0;
wire [15:0] PE151_out1;
wire [15:0] PE151_out2;
wire [15:0] PE151_out3;

wire [15:0] PE152_out0;
wire [15:0] PE152_out1;
wire [15:0] PE152_out2;
wire [15:0] PE152_out3;

wire [15:0] PE153_out0;
wire [15:0] PE153_out1;
wire [15:0] PE153_out2;
wire [15:0] PE153_out3;

wire [15:0] PE154_out0;
wire [15:0] PE154_out1;
wire [15:0] PE154_out2;
wire [15:0] PE154_out3;

wire [15:0] PE155_out0;
wire [15:0] PE155_out1;
wire [15:0] PE155_out2;
wire [15:0] PE155_out3;

wire [15:0] PE156_out0;
wire [15:0] PE156_out1;
wire [15:0] PE156_out2;
wire [15:0] PE156_out3;

wire [15:0] PE157_out0;
wire [15:0] PE157_out1;
wire [15:0] PE157_out2;
wire [15:0] PE157_out3;



PE PE00(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE07_out2),
     .PE_in1(PE150_out3),
     .PE_in2(PE01_out0),
     .PE_in3(PE10_out1),

     .PE_out0(PE00_out0),
     .PE_out1(PE00_out1),
     .PE_out2(PE00_out2),
     .PE_out3(PE00_out3)
       );

PE PE01(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE00_out2),
     .PE_in1(PE151_out3),
     .PE_in2(PE02_out0),
     .PE_in3(PE11_out1),

     .PE_out0(PE01_out0),
     .PE_out1(PE01_out1),
     .PE_out2(PE01_out2),
     .PE_out3(PE01_out3)
       );

PE PE02(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE01_out2),
     .PE_in1(PE152_out3),
     .PE_in2(PE03_out0),
     .PE_in3(PE12_out1),

     .PE_out0(PE02_out0),
     .PE_out1(PE02_out1),
     .PE_out2(PE02_out2),
     .PE_out3(PE02_out3)
       );

PE PE03(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE02_out2),
     .PE_in1(PE153_out3),
     .PE_in2(PE04_out0),
     .PE_in3(PE13_out1),

     .PE_out0(PE03_out0),
     .PE_out1(PE03_out1),
     .PE_out2(PE03_out2),
     .PE_out3(PE03_out3)
       );

PE PE04(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE03_out2),
     .PE_in1(PE154_out3),
     .PE_in2(PE05_out0),
     .PE_in3(PE14_out1),

     .PE_out0(PE04_out0),
     .PE_out1(PE04_out1),
     .PE_out2(PE04_out2),
     .PE_out3(PE04_out3)
       );

PE PE05(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE04_out2),
     .PE_in1(PE155_out3),
     .PE_in2(PE06_out0),
     .PE_in3(PE15_out1),

     .PE_out0(PE05_out0),
     .PE_out1(PE05_out1),
     .PE_out2(PE05_out2),
     .PE_out3(PE05_out3)
       );

PE PE06(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE05_out2),
     .PE_in1(PE156_out3),
     .PE_in2(PE07_out0),
     .PE_in3(PE16_out1),

     .PE_out0(PE06_out0),
     .PE_out1(PE06_out1),
     .PE_out2(PE06_out2),
     .PE_out3(PE06_out3)
       );

PE PE07(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE06_out2),
     .PE_in1(PE157_out3),
     .PE_in2(PE00_out0),
     .PE_in3(PE17_out1),

     .PE_out0(PE07_out0),
     .PE_out1(PE07_out1),
     .PE_out2(PE07_out2),
     .PE_out3(PE07_out3)
       );


PE PE10(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE17_out2),
     .PE_in1(PE00_out3),
     .PE_in2(PE11_out0),
     .PE_in3(PE20_out1),

     .PE_out0(PE10_out0),
     .PE_out1(PE10_out1),
     .PE_out2(PE10_out2),
     .PE_out3(PE10_out3)
       );

PE PE11(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE10_out2),
     .PE_in1(PE01_out3),
     .PE_in2(PE12_out0),
     .PE_in3(PE21_out1),

     .PE_out0(PE11_out0),
     .PE_out1(PE11_out1),
     .PE_out2(PE11_out2),
     .PE_out3(PE11_out3)
       );

PE PE12(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE11_out2),
     .PE_in1(PE02_out3),
     .PE_in2(PE13_out0),
     .PE_in3(PE22_out1),

     .PE_out0(PE12_out0),
     .PE_out1(PE12_out1),
     .PE_out2(PE12_out2),
     .PE_out3(PE12_out3)
       );

PE PE13(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE12_out2),
     .PE_in1(PE03_out3),
     .PE_in2(PE14_out0),
     .PE_in3(PE23_out1),

     .PE_out0(PE13_out0),
     .PE_out1(PE13_out1),
     .PE_out2(PE13_out2),
     .PE_out3(PE13_out3)
       );

PE PE14(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE13_out2),
     .PE_in1(PE04_out3),
     .PE_in2(PE15_out0),
     .PE_in3(PE24_out1),

     .PE_out0(PE14_out0),
     .PE_out1(PE14_out1),
     .PE_out2(PE14_out2),
     .PE_out3(PE14_out3)
       );

PE PE15(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE14_out2),
     .PE_in1(PE05_out3),
     .PE_in2(PE16_out0),
     .PE_in3(PE25_out1),

     .PE_out0(PE15_out0),
     .PE_out1(PE15_out1),
     .PE_out2(PE15_out2),
     .PE_out3(PE15_out3)
       );

PE PE16(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE15_out2),
     .PE_in1(PE06_out3),
     .PE_in2(PE17_out0),
     .PE_in3(PE26_out1),

     .PE_out0(PE16_out0),
     .PE_out1(PE16_out1),
     .PE_out2(PE16_out2),
     .PE_out3(PE16_out3)
       );

PE PE17(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE16_out2),
     .PE_in1(PE07_out3),
     .PE_in2(PE10_out0),
     .PE_in3(PE27_out1),

     .PE_out0(PE17_out0),
     .PE_out1(PE17_out1),
     .PE_out2(PE17_out2),
     .PE_out3(PE17_out3)
       );


PE PE20(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE27_out2),
     .PE_in1(PE10_out3),
     .PE_in2(PE21_out0),
     .PE_in3(PE30_out1),

     .PE_out0(PE20_out0),
     .PE_out1(PE20_out1),
     .PE_out2(PE20_out2),
     .PE_out3(PE20_out3)
       );

PE PE21(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE20_out2),
     .PE_in1(PE11_out3),
     .PE_in2(PE22_out0),
     .PE_in3(PE31_out1),

     .PE_out0(PE21_out0),
     .PE_out1(PE21_out1),
     .PE_out2(PE21_out2),
     .PE_out3(PE21_out3)
       );

PE PE22(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE21_out2),
     .PE_in1(PE12_out3),
     .PE_in2(PE23_out0),
     .PE_in3(PE32_out1),

     .PE_out0(PE22_out0),
     .PE_out1(PE22_out1),
     .PE_out2(PE22_out2),
     .PE_out3(PE22_out3)
       );

PE PE23(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE22_out2),
     .PE_in1(PE13_out3),
     .PE_in2(PE24_out0),
     .PE_in3(PE33_out1),

     .PE_out0(PE23_out0),
     .PE_out1(PE23_out1),
     .PE_out2(PE23_out2),
     .PE_out3(PE23_out3)
       );

PE PE24(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE23_out2),
     .PE_in1(PE14_out3),
     .PE_in2(PE25_out0),
     .PE_in3(PE34_out1),

     .PE_out0(PE24_out0),
     .PE_out1(PE24_out1),
     .PE_out2(PE24_out2),
     .PE_out3(PE24_out3)
       );

PE PE25(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE24_out2),
     .PE_in1(PE15_out3),
     .PE_in2(PE26_out0),
     .PE_in3(PE35_out1),

     .PE_out0(PE25_out0),
     .PE_out1(PE25_out1),
     .PE_out2(PE25_out2),
     .PE_out3(PE25_out3)
       );

PE PE26(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE25_out2),
     .PE_in1(PE16_out3),
     .PE_in2(PE27_out0),
     .PE_in3(PE36_out1),

     .PE_out0(PE26_out0),
     .PE_out1(PE26_out1),
     .PE_out2(PE26_out2),
     .PE_out3(PE26_out3)
       );

PE PE27(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE26_out2),
     .PE_in1(PE17_out3),
     .PE_in2(PE20_out0),
     .PE_in3(PE37_out1),

     .PE_out0(PE27_out0),
     .PE_out1(PE27_out1),
     .PE_out2(PE27_out2),
     .PE_out3(PE27_out3)
       );


PE PE30(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE37_out2),
     .PE_in1(PE20_out3),
     .PE_in2(PE31_out0),
     .PE_in3(PE40_out1),

     .PE_out0(PE30_out0),
     .PE_out1(PE30_out1),
     .PE_out2(PE30_out2),
     .PE_out3(PE30_out3)
       );

PE PE31(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE30_out2),
     .PE_in1(PE21_out3),
     .PE_in2(PE32_out0),
     .PE_in3(PE41_out1),

     .PE_out0(PE31_out0),
     .PE_out1(PE31_out1),
     .PE_out2(PE31_out2),
     .PE_out3(PE31_out3)
       );

PE PE32(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE31_out2),
     .PE_in1(PE22_out3),
     .PE_in2(PE33_out0),
     .PE_in3(PE42_out1),

     .PE_out0(PE32_out0),
     .PE_out1(PE32_out1),
     .PE_out2(PE32_out2),
     .PE_out3(PE32_out3)
       );

PE PE33(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE32_out2),
     .PE_in1(PE23_out3),
     .PE_in2(PE34_out0),
     .PE_in3(PE43_out1),

     .PE_out0(PE33_out0),
     .PE_out1(PE33_out1),
     .PE_out2(PE33_out2),
     .PE_out3(PE33_out3)
       );

PE PE34(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE33_out2),
     .PE_in1(PE24_out3),
     .PE_in2(PE35_out0),
     .PE_in3(PE44_out1),

     .PE_out0(PE34_out0),
     .PE_out1(PE34_out1),
     .PE_out2(PE34_out2),
     .PE_out3(PE34_out3)
       );

PE PE35(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE34_out2),
     .PE_in1(PE25_out3),
     .PE_in2(PE36_out0),
     .PE_in3(PE45_out1),

     .PE_out0(PE35_out0),
     .PE_out1(PE35_out1),
     .PE_out2(PE35_out2),
     .PE_out3(PE35_out3)
       );

PE PE36(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE35_out2),
     .PE_in1(PE26_out3),
     .PE_in2(PE37_out0),
     .PE_in3(PE46_out1),

     .PE_out0(PE36_out0),
     .PE_out1(PE36_out1),
     .PE_out2(PE36_out2),
     .PE_out3(PE36_out3)
       );

PE PE37(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE36_out2),
     .PE_in1(PE27_out3),
     .PE_in2(PE30_out0),
     .PE_in3(PE47_out1),

     .PE_out0(PE37_out0),
     .PE_out1(PE37_out1),
     .PE_out2(PE37_out2),
     .PE_out3(PE37_out3)
       );


PE PE40(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE47_out2),
     .PE_in1(PE30_out3),
     .PE_in2(PE41_out0),
     .PE_in3(PE50_out1),

     .PE_out0(PE40_out0),
     .PE_out1(PE40_out1),
     .PE_out2(PE40_out2),
     .PE_out3(PE40_out3)
       );

PE PE41(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE40_out2),
     .PE_in1(PE31_out3),
     .PE_in2(PE42_out0),
     .PE_in3(PE51_out1),

     .PE_out0(PE41_out0),
     .PE_out1(PE41_out1),
     .PE_out2(PE41_out2),
     .PE_out3(PE41_out3)
       );

PE PE42(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE41_out2),
     .PE_in1(PE32_out3),
     .PE_in2(PE43_out0),
     .PE_in3(PE52_out1),

     .PE_out0(PE42_out0),
     .PE_out1(PE42_out1),
     .PE_out2(PE42_out2),
     .PE_out3(PE42_out3)
       );

PE PE43(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE42_out2),
     .PE_in1(PE33_out3),
     .PE_in2(PE44_out0),
     .PE_in3(PE53_out1),

     .PE_out0(PE43_out0),
     .PE_out1(PE43_out1),
     .PE_out2(PE43_out2),
     .PE_out3(PE43_out3)
       );

PE PE44(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE43_out2),
     .PE_in1(PE34_out3),
     .PE_in2(PE45_out0),
     .PE_in3(PE54_out1),

     .PE_out0(PE44_out0),
     .PE_out1(PE44_out1),
     .PE_out2(PE44_out2),
     .PE_out3(PE44_out3)
       );

PE PE45(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE44_out2),
     .PE_in1(PE35_out3),
     .PE_in2(PE46_out0),
     .PE_in3(PE55_out1),

     .PE_out0(PE45_out0),
     .PE_out1(PE45_out1),
     .PE_out2(PE45_out2),
     .PE_out3(PE45_out3)
       );

PE PE46(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE45_out2),
     .PE_in1(PE36_out3),
     .PE_in2(PE47_out0),
     .PE_in3(PE56_out1),

     .PE_out0(PE46_out0),
     .PE_out1(PE46_out1),
     .PE_out2(PE46_out2),
     .PE_out3(PE46_out3)
       );

PE PE47(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE46_out2),
     .PE_in1(PE37_out3),
     .PE_in2(PE40_out0),
     .PE_in3(PE57_out1),

     .PE_out0(PE47_out0),
     .PE_out1(PE47_out1),
     .PE_out2(PE47_out2),
     .PE_out3(PE47_out3)
       );


PE PE50(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE57_out2),
     .PE_in1(PE40_out3),
     .PE_in2(PE51_out0),
     .PE_in3(PE60_out1),

     .PE_out0(PE50_out0),
     .PE_out1(PE50_out1),
     .PE_out2(PE50_out2),
     .PE_out3(PE50_out3)
       );

PE PE51(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE50_out2),
     .PE_in1(PE41_out3),
     .PE_in2(PE52_out0),
     .PE_in3(PE61_out1),

     .PE_out0(PE51_out0),
     .PE_out1(PE51_out1),
     .PE_out2(PE51_out2),
     .PE_out3(PE51_out3)
       );

PE PE52(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE51_out2),
     .PE_in1(PE42_out3),
     .PE_in2(PE53_out0),
     .PE_in3(PE62_out1),

     .PE_out0(PE52_out0),
     .PE_out1(PE52_out1),
     .PE_out2(PE52_out2),
     .PE_out3(PE52_out3)
       );

PE PE53(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE52_out2),
     .PE_in1(PE43_out3),
     .PE_in2(PE54_out0),
     .PE_in3(PE63_out1),

     .PE_out0(PE53_out0),
     .PE_out1(PE53_out1),
     .PE_out2(PE53_out2),
     .PE_out3(PE53_out3)
       );

PE PE54(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE53_out2),
     .PE_in1(PE44_out3),
     .PE_in2(PE55_out0),
     .PE_in3(PE64_out1),

     .PE_out0(PE54_out0),
     .PE_out1(PE54_out1),
     .PE_out2(PE54_out2),
     .PE_out3(PE54_out3)
       );

PE PE55(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE54_out2),
     .PE_in1(PE45_out3),
     .PE_in2(PE56_out0),
     .PE_in3(PE65_out1),

     .PE_out0(PE55_out0),
     .PE_out1(PE55_out1),
     .PE_out2(PE55_out2),
     .PE_out3(PE55_out3)
       );

PE PE56(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE55_out2),
     .PE_in1(PE46_out3),
     .PE_in2(PE57_out0),
     .PE_in3(PE66_out1),

     .PE_out0(PE56_out0),
     .PE_out1(PE56_out1),
     .PE_out2(PE56_out2),
     .PE_out3(PE56_out3)
       );

PE PE57(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE56_out2),
     .PE_in1(PE47_out3),
     .PE_in2(PE50_out0),
     .PE_in3(PE67_out1),

     .PE_out0(PE57_out0),
     .PE_out1(PE57_out1),
     .PE_out2(PE57_out2),
     .PE_out3(PE57_out3)
       );


PE PE60(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE67_out2),
     .PE_in1(PE50_out3),
     .PE_in2(PE61_out0),
     .PE_in3(PE70_out1),

     .PE_out0(PE60_out0),
     .PE_out1(PE60_out1),
     .PE_out2(PE60_out2),
     .PE_out3(PE60_out3)
       );

PE PE61(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE60_out2),
     .PE_in1(PE51_out3),
     .PE_in2(PE62_out0),
     .PE_in3(PE71_out1),

     .PE_out0(PE61_out0),
     .PE_out1(PE61_out1),
     .PE_out2(PE61_out2),
     .PE_out3(PE61_out3)
       );

PE PE62(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE61_out2),
     .PE_in1(PE52_out3),
     .PE_in2(PE63_out0),
     .PE_in3(PE72_out1),

     .PE_out0(PE62_out0),
     .PE_out1(PE62_out1),
     .PE_out2(PE62_out2),
     .PE_out3(PE62_out3)
       );

PE PE63(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE62_out2),
     .PE_in1(PE53_out3),
     .PE_in2(PE64_out0),
     .PE_in3(PE73_out1),

     .PE_out0(PE63_out0),
     .PE_out1(PE63_out1),
     .PE_out2(PE63_out2),
     .PE_out3(PE63_out3)
       );

PE PE64(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE63_out2),
     .PE_in1(PE54_out3),
     .PE_in2(PE65_out0),
     .PE_in3(PE74_out1),

     .PE_out0(PE64_out0),
     .PE_out1(PE64_out1),
     .PE_out2(PE64_out2),
     .PE_out3(PE64_out3)
       );

PE PE65(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE64_out2),
     .PE_in1(PE55_out3),
     .PE_in2(PE66_out0),
     .PE_in3(PE75_out1),

     .PE_out0(PE65_out0),
     .PE_out1(PE65_out1),
     .PE_out2(PE65_out2),
     .PE_out3(PE65_out3)
       );

PE PE66(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE65_out2),
     .PE_in1(PE56_out3),
     .PE_in2(PE67_out0),
     .PE_in3(PE76_out1),

     .PE_out0(PE66_out0),
     .PE_out1(PE66_out1),
     .PE_out2(PE66_out2),
     .PE_out3(PE66_out3)
       );

PE PE67(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE66_out2),
     .PE_in1(PE57_out3),
     .PE_in2(PE60_out0),
     .PE_in3(PE77_out1),

     .PE_out0(PE67_out0),
     .PE_out1(PE67_out1),
     .PE_out2(PE67_out2),
     .PE_out3(PE67_out3)
       );


PE PE70(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE77_out2),
     .PE_in1(PE60_out3),
     .PE_in2(PE71_out0),
     .PE_in3(PE80_out1),

     .PE_out0(PE70_out0),
     .PE_out1(PE70_out1),
     .PE_out2(PE70_out2),
     .PE_out3(PE70_out3)
       );

PE PE71(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE70_out2),
     .PE_in1(PE61_out3),
     .PE_in2(PE72_out0),
     .PE_in3(PE81_out1),

     .PE_out0(PE71_out0),
     .PE_out1(PE71_out1),
     .PE_out2(PE71_out2),
     .PE_out3(PE71_out3)
       );

PE PE72(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE71_out2),
     .PE_in1(PE62_out3),
     .PE_in2(PE73_out0),
     .PE_in3(PE82_out1),

     .PE_out0(PE72_out0),
     .PE_out1(PE72_out1),
     .PE_out2(PE72_out2),
     .PE_out3(PE72_out3)
       );

PE PE73(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE72_out2),
     .PE_in1(PE63_out3),
     .PE_in2(PE74_out0),
     .PE_in3(PE83_out1),

     .PE_out0(PE73_out0),
     .PE_out1(PE73_out1),
     .PE_out2(PE73_out2),
     .PE_out3(PE73_out3)
       );

PE PE74(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE73_out2),
     .PE_in1(PE64_out3),
     .PE_in2(PE75_out0),
     .PE_in3(PE84_out1),

     .PE_out0(PE74_out0),
     .PE_out1(PE74_out1),
     .PE_out2(PE74_out2),
     .PE_out3(PE74_out3)
       );

PE PE75(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE74_out2),
     .PE_in1(PE65_out3),
     .PE_in2(PE76_out0),
     .PE_in3(PE85_out1),

     .PE_out0(PE75_out0),
     .PE_out1(PE75_out1),
     .PE_out2(PE75_out2),
     .PE_out3(PE75_out3)
       );

PE PE76(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE75_out2),
     .PE_in1(PE66_out3),
     .PE_in2(PE77_out0),
     .PE_in3(PE86_out1),

     .PE_out0(PE76_out0),
     .PE_out1(PE76_out1),
     .PE_out2(PE76_out2),
     .PE_out3(PE76_out3)
       );

PE PE77(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE76_out2),
     .PE_in1(PE67_out3),
     .PE_in2(PE70_out0),
     .PE_in3(PE87_out1),

     .PE_out0(PE77_out0),
     .PE_out1(PE77_out1),
     .PE_out2(PE77_out2),
     .PE_out3(PE77_out3)
       );


PE PE80(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE87_out2),
     .PE_in1(PE70_out3),
     .PE_in2(PE81_out0),
     .PE_in3(PE90_out1),

     .PE_out0(PE80_out0),
     .PE_out1(PE80_out1),
     .PE_out2(PE80_out2),
     .PE_out3(PE80_out3)
       );

PE PE81(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE80_out2),
     .PE_in1(PE71_out3),
     .PE_in2(PE82_out0),
     .PE_in3(PE91_out1),

     .PE_out0(PE81_out0),
     .PE_out1(PE81_out1),
     .PE_out2(PE81_out2),
     .PE_out3(PE81_out3)
       );

PE PE82(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE81_out2),
     .PE_in1(PE72_out3),
     .PE_in2(PE83_out0),
     .PE_in3(PE92_out1),

     .PE_out0(PE82_out0),
     .PE_out1(PE82_out1),
     .PE_out2(PE82_out2),
     .PE_out3(PE82_out3)
       );

PE PE83(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE82_out2),
     .PE_in1(PE73_out3),
     .PE_in2(PE84_out0),
     .PE_in3(PE93_out1),

     .PE_out0(PE83_out0),
     .PE_out1(PE83_out1),
     .PE_out2(PE83_out2),
     .PE_out3(PE83_out3)
       );

PE PE84(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE83_out2),
     .PE_in1(PE74_out3),
     .PE_in2(PE85_out0),
     .PE_in3(PE94_out1),

     .PE_out0(PE84_out0),
     .PE_out1(PE84_out1),
     .PE_out2(PE84_out2),
     .PE_out3(PE84_out3)
       );

PE PE85(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE84_out2),
     .PE_in1(PE75_out3),
     .PE_in2(PE86_out0),
     .PE_in3(PE95_out1),

     .PE_out0(PE85_out0),
     .PE_out1(PE85_out1),
     .PE_out2(PE85_out2),
     .PE_out3(PE85_out3)
       );

PE PE86(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE85_out2),
     .PE_in1(PE76_out3),
     .PE_in2(PE87_out0),
     .PE_in3(PE96_out1),

     .PE_out0(PE86_out0),
     .PE_out1(PE86_out1),
     .PE_out2(PE86_out2),
     .PE_out3(PE86_out3)
       );

PE PE87(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE86_out2),
     .PE_in1(PE77_out3),
     .PE_in2(PE80_out0),
     .PE_in3(PE97_out1),

     .PE_out0(PE87_out0),
     .PE_out1(PE87_out1),
     .PE_out2(PE87_out2),
     .PE_out3(PE87_out3)
       );


PE PE90(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE97_out2),
     .PE_in1(PE80_out3),
     .PE_in2(PE91_out0),
     .PE_in3(PE100_out1),

     .PE_out0(PE90_out0),
     .PE_out1(PE90_out1),
     .PE_out2(PE90_out2),
     .PE_out3(PE90_out3)
       );

PE PE91(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE90_out2),
     .PE_in1(PE81_out3),
     .PE_in2(PE92_out0),
     .PE_in3(PE101_out1),

     .PE_out0(PE91_out0),
     .PE_out1(PE91_out1),
     .PE_out2(PE91_out2),
     .PE_out3(PE91_out3)
       );

PE PE92(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE91_out2),
     .PE_in1(PE82_out3),
     .PE_in2(PE93_out0),
     .PE_in3(PE102_out1),

     .PE_out0(PE92_out0),
     .PE_out1(PE92_out1),
     .PE_out2(PE92_out2),
     .PE_out3(PE92_out3)
       );

PE PE93(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE92_out2),
     .PE_in1(PE83_out3),
     .PE_in2(PE94_out0),
     .PE_in3(PE103_out1),

     .PE_out0(PE93_out0),
     .PE_out1(PE93_out1),
     .PE_out2(PE93_out2),
     .PE_out3(PE93_out3)
       );

PE PE94(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE93_out2),
     .PE_in1(PE84_out3),
     .PE_in2(PE95_out0),
     .PE_in3(PE104_out1),

     .PE_out0(PE94_out0),
     .PE_out1(PE94_out1),
     .PE_out2(PE94_out2),
     .PE_out3(PE94_out3)
       );

PE PE95(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE94_out2),
     .PE_in1(PE85_out3),
     .PE_in2(PE96_out0),
     .PE_in3(PE105_out1),

     .PE_out0(PE95_out0),
     .PE_out1(PE95_out1),
     .PE_out2(PE95_out2),
     .PE_out3(PE95_out3)
       );

PE PE96(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE95_out2),
     .PE_in1(PE86_out3),
     .PE_in2(PE97_out0),
     .PE_in3(PE106_out1),

     .PE_out0(PE96_out0),
     .PE_out1(PE96_out1),
     .PE_out2(PE96_out2),
     .PE_out3(PE96_out3)
       );

PE PE97(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE96_out2),
     .PE_in1(PE87_out3),
     .PE_in2(PE90_out0),
     .PE_in3(PE107_out1),

     .PE_out0(PE97_out0),
     .PE_out1(PE97_out1),
     .PE_out2(PE97_out2),
     .PE_out3(PE97_out3)
       );


PE PE100(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE107_out2),
     .PE_in1(PE90_out3),
     .PE_in2(PE101_out0),
     .PE_in3(PE110_out1),

     .PE_out0(PE100_out0),
     .PE_out1(PE100_out1),
     .PE_out2(PE100_out2),
     .PE_out3(PE100_out3)
       );

PE PE101(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE100_out2),
     .PE_in1(PE91_out3),
     .PE_in2(PE102_out0),
     .PE_in3(PE111_out1),

     .PE_out0(PE101_out0),
     .PE_out1(PE101_out1),
     .PE_out2(PE101_out2),
     .PE_out3(PE101_out3)
       );

PE PE102(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE101_out2),
     .PE_in1(PE92_out3),
     .PE_in2(PE103_out0),
     .PE_in3(PE112_out1),

     .PE_out0(PE102_out0),
     .PE_out1(PE102_out1),
     .PE_out2(PE102_out2),
     .PE_out3(PE102_out3)
       );

PE PE103(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE102_out2),
     .PE_in1(PE93_out3),
     .PE_in2(PE104_out0),
     .PE_in3(PE113_out1),

     .PE_out0(PE103_out0),
     .PE_out1(PE103_out1),
     .PE_out2(PE103_out2),
     .PE_out3(PE103_out3)
       );

PE PE104(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE103_out2),
     .PE_in1(PE94_out3),
     .PE_in2(PE105_out0),
     .PE_in3(PE114_out1),

     .PE_out0(PE104_out0),
     .PE_out1(PE104_out1),
     .PE_out2(PE104_out2),
     .PE_out3(PE104_out3)
       );

PE PE105(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE104_out2),
     .PE_in1(PE95_out3),
     .PE_in2(PE106_out0),
     .PE_in3(PE115_out1),

     .PE_out0(PE105_out0),
     .PE_out1(PE105_out1),
     .PE_out2(PE105_out2),
     .PE_out3(PE105_out3)
       );

PE PE106(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE105_out2),
     .PE_in1(PE96_out3),
     .PE_in2(PE107_out0),
     .PE_in3(PE116_out1),

     .PE_out0(PE106_out0),
     .PE_out1(PE106_out1),
     .PE_out2(PE106_out2),
     .PE_out3(PE106_out3)
       );

PE PE107(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE106_out2),
     .PE_in1(PE97_out3),
     .PE_in2(PE100_out0),
     .PE_in3(PE117_out1),

     .PE_out0(PE107_out0),
     .PE_out1(PE107_out1),
     .PE_out2(PE107_out2),
     .PE_out3(PE107_out3)
       );


PE PE110(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE117_out2),
     .PE_in1(PE100_out3),
     .PE_in2(PE111_out0),
     .PE_in3(PE120_out1),

     .PE_out0(PE110_out0),
     .PE_out1(PE110_out1),
     .PE_out2(PE110_out2),
     .PE_out3(PE110_out3)
       );

PE PE111(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE110_out2),
     .PE_in1(PE101_out3),
     .PE_in2(PE112_out0),
     .PE_in3(PE121_out1),

     .PE_out0(PE111_out0),
     .PE_out1(PE111_out1),
     .PE_out2(PE111_out2),
     .PE_out3(PE111_out3)
       );

PE PE112(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE111_out2),
     .PE_in1(PE102_out3),
     .PE_in2(PE113_out0),
     .PE_in3(PE122_out1),

     .PE_out0(PE112_out0),
     .PE_out1(PE112_out1),
     .PE_out2(PE112_out2),
     .PE_out3(PE112_out3)
       );

PE PE113(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE112_out2),
     .PE_in1(PE103_out3),
     .PE_in2(PE114_out0),
     .PE_in3(PE123_out1),

     .PE_out0(PE113_out0),
     .PE_out1(PE113_out1),
     .PE_out2(PE113_out2),
     .PE_out3(PE113_out3)
       );

PE PE114(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE113_out2),
     .PE_in1(PE104_out3),
     .PE_in2(PE115_out0),
     .PE_in3(PE124_out1),

     .PE_out0(PE114_out0),
     .PE_out1(PE114_out1),
     .PE_out2(PE114_out2),
     .PE_out3(PE114_out3)
       );

PE PE115(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE114_out2),
     .PE_in1(PE105_out3),
     .PE_in2(PE116_out0),
     .PE_in3(PE125_out1),

     .PE_out0(PE115_out0),
     .PE_out1(PE115_out1),
     .PE_out2(PE115_out2),
     .PE_out3(PE115_out3)
       );

PE PE116(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE115_out2),
     .PE_in1(PE106_out3),
     .PE_in2(PE117_out0),
     .PE_in3(PE126_out1),

     .PE_out0(PE116_out0),
     .PE_out1(PE116_out1),
     .PE_out2(PE116_out2),
     .PE_out3(PE116_out3)
       );

PE PE117(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE116_out2),
     .PE_in1(PE107_out3),
     .PE_in2(PE110_out0),
     .PE_in3(PE127_out1),

     .PE_out0(PE117_out0),
     .PE_out1(PE117_out1),
     .PE_out2(PE117_out2),
     .PE_out3(PE117_out3)
       );


PE PE120(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE127_out2),
     .PE_in1(PE110_out3),
     .PE_in2(PE121_out0),
     .PE_in3(PE130_out1),

     .PE_out0(PE120_out0),
     .PE_out1(PE120_out1),
     .PE_out2(PE120_out2),
     .PE_out3(PE120_out3)
       );

PE PE121(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE120_out2),
     .PE_in1(PE111_out3),
     .PE_in2(PE122_out0),
     .PE_in3(PE131_out1),

     .PE_out0(PE121_out0),
     .PE_out1(PE121_out1),
     .PE_out2(PE121_out2),
     .PE_out3(PE121_out3)
       );

PE PE122(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE121_out2),
     .PE_in1(PE112_out3),
     .PE_in2(PE123_out0),
     .PE_in3(PE132_out1),

     .PE_out0(PE122_out0),
     .PE_out1(PE122_out1),
     .PE_out2(PE122_out2),
     .PE_out3(PE122_out3)
       );

PE PE123(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE122_out2),
     .PE_in1(PE113_out3),
     .PE_in2(PE124_out0),
     .PE_in3(PE133_out1),

     .PE_out0(PE123_out0),
     .PE_out1(PE123_out1),
     .PE_out2(PE123_out2),
     .PE_out3(PE123_out3)
       );

PE PE124(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE123_out2),
     .PE_in1(PE114_out3),
     .PE_in2(PE125_out0),
     .PE_in3(PE134_out1),

     .PE_out0(PE124_out0),
     .PE_out1(PE124_out1),
     .PE_out2(PE124_out2),
     .PE_out3(PE124_out3)
       );

PE PE125(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE124_out2),
     .PE_in1(PE115_out3),
     .PE_in2(PE126_out0),
     .PE_in3(PE135_out1),

     .PE_out0(PE125_out0),
     .PE_out1(PE125_out1),
     .PE_out2(PE125_out2),
     .PE_out3(PE125_out3)
       );

PE PE126(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE125_out2),
     .PE_in1(PE116_out3),
     .PE_in2(PE127_out0),
     .PE_in3(PE136_out1),

     .PE_out0(PE126_out0),
     .PE_out1(PE126_out1),
     .PE_out2(PE126_out2),
     .PE_out3(PE126_out3)
       );

PE PE127(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE126_out2),
     .PE_in1(PE117_out3),
     .PE_in2(PE120_out0),
     .PE_in3(PE137_out1),

     .PE_out0(PE127_out0),
     .PE_out1(PE127_out1),
     .PE_out2(PE127_out2),
     .PE_out3(PE127_out3)
       );


PE PE130(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE137_out2),
     .PE_in1(PE120_out3),
     .PE_in2(PE131_out0),
     .PE_in3(PE140_out1),

     .PE_out0(PE130_out0),
     .PE_out1(PE130_out1),
     .PE_out2(PE130_out2),
     .PE_out3(PE130_out3)
       );

PE PE131(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE130_out2),
     .PE_in1(PE121_out3),
     .PE_in2(PE132_out0),
     .PE_in3(PE141_out1),

     .PE_out0(PE131_out0),
     .PE_out1(PE131_out1),
     .PE_out2(PE131_out2),
     .PE_out3(PE131_out3)
       );

PE PE132(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE131_out2),
     .PE_in1(PE122_out3),
     .PE_in2(PE133_out0),
     .PE_in3(PE142_out1),

     .PE_out0(PE132_out0),
     .PE_out1(PE132_out1),
     .PE_out2(PE132_out2),
     .PE_out3(PE132_out3)
       );

PE PE133(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE132_out2),
     .PE_in1(PE123_out3),
     .PE_in2(PE134_out0),
     .PE_in3(PE143_out1),

     .PE_out0(PE133_out0),
     .PE_out1(PE133_out1),
     .PE_out2(PE133_out2),
     .PE_out3(PE133_out3)
       );

PE PE134(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE133_out2),
     .PE_in1(PE124_out3),
     .PE_in2(PE135_out0),
     .PE_in3(PE144_out1),

     .PE_out0(PE134_out0),
     .PE_out1(PE134_out1),
     .PE_out2(PE134_out2),
     .PE_out3(PE134_out3)
       );

PE PE135(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE134_out2),
     .PE_in1(PE125_out3),
     .PE_in2(PE136_out0),
     .PE_in3(PE145_out1),

     .PE_out0(PE135_out0),
     .PE_out1(PE135_out1),
     .PE_out2(PE135_out2),
     .PE_out3(PE135_out3)
       );

PE PE136(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE135_out2),
     .PE_in1(PE126_out3),
     .PE_in2(PE137_out0),
     .PE_in3(PE146_out1),

     .PE_out0(PE136_out0),
     .PE_out1(PE136_out1),
     .PE_out2(PE136_out2),
     .PE_out3(PE136_out3)
       );

PE PE137(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE136_out2),
     .PE_in1(PE127_out3),
     .PE_in2(PE130_out0),
     .PE_in3(PE147_out1),

     .PE_out0(PE137_out0),
     .PE_out1(PE137_out1),
     .PE_out2(PE137_out2),
     .PE_out3(PE137_out3)
       );


PE PE140(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE147_out2),
     .PE_in1(PE130_out3),
     .PE_in2(PE141_out0),
     .PE_in3(PE150_out1),

     .PE_out0(PE140_out0),
     .PE_out1(PE140_out1),
     .PE_out2(PE140_out2),
     .PE_out3(PE140_out3)
       );

PE PE141(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE140_out2),
     .PE_in1(PE131_out3),
     .PE_in2(PE142_out0),
     .PE_in3(PE151_out1),

     .PE_out0(PE141_out0),
     .PE_out1(PE141_out1),
     .PE_out2(PE141_out2),
     .PE_out3(PE141_out3)
       );

PE PE142(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE141_out2),
     .PE_in1(PE132_out3),
     .PE_in2(PE143_out0),
     .PE_in3(PE152_out1),

     .PE_out0(PE142_out0),
     .PE_out1(PE142_out1),
     .PE_out2(PE142_out2),
     .PE_out3(PE142_out3)
       );

PE PE143(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE142_out2),
     .PE_in1(PE133_out3),
     .PE_in2(PE144_out0),
     .PE_in3(PE153_out1),

     .PE_out0(PE143_out0),
     .PE_out1(PE143_out1),
     .PE_out2(PE143_out2),
     .PE_out3(PE143_out3)
       );

PE PE144(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE143_out2),
     .PE_in1(PE134_out3),
     .PE_in2(PE145_out0),
     .PE_in3(PE154_out1),

     .PE_out0(PE144_out0),
     .PE_out1(PE144_out1),
     .PE_out2(PE144_out2),
     .PE_out3(PE144_out3)
       );

PE PE145(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE144_out2),
     .PE_in1(PE135_out3),
     .PE_in2(PE146_out0),
     .PE_in3(PE155_out1),

     .PE_out0(PE145_out0),
     .PE_out1(PE145_out1),
     .PE_out2(PE145_out2),
     .PE_out3(PE145_out3)
       );

PE PE146(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE145_out2),
     .PE_in1(PE136_out3),
     .PE_in2(PE147_out0),
     .PE_in3(PE156_out1),

     .PE_out0(PE146_out0),
     .PE_out1(PE146_out1),
     .PE_out2(PE146_out2),
     .PE_out3(PE146_out3)
       );

PE PE147(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE146_out2),
     .PE_in1(PE137_out3),
     .PE_in2(PE140_out0),
     .PE_in3(PE157_out1),

     .PE_out0(PE147_out0),
     .PE_out1(PE147_out1),
     .PE_out2(PE147_out2),
     .PE_out3(PE147_out3)
       );


PE PE150(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE157_out2),
     .PE_in1(PE140_out3),
     .PE_in2(PE151_out0),
     .PE_in3(PE00_out1),

     .PE_out0(PE150_out0),
     .PE_out1(PE150_out1),
     .PE_out2(PE150_out2),
     .PE_out3(PE150_out3)
       );

PE PE151(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE150_out2),
     .PE_in1(PE141_out3),
     .PE_in2(PE152_out0),
     .PE_in3(PE01_out1),

     .PE_out0(PE151_out0),
     .PE_out1(PE151_out1),
     .PE_out2(PE151_out2),
     .PE_out3(PE151_out3)
       );

PE PE152(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE151_out2),
     .PE_in1(PE142_out3),
     .PE_in2(PE153_out0),
     .PE_in3(PE02_out1),

     .PE_out0(PE152_out0),
     .PE_out1(PE152_out1),
     .PE_out2(PE152_out2),
     .PE_out3(PE152_out3)
       );

PE PE153(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE152_out2),
     .PE_in1(PE143_out3),
     .PE_in2(PE154_out0),
     .PE_in3(PE03_out1),

     .PE_out0(PE153_out0),
     .PE_out1(PE153_out1),
     .PE_out2(PE153_out2),
     .PE_out3(PE153_out3)
       );

PE PE154(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE153_out2),
     .PE_in1(PE144_out3),
     .PE_in2(PE155_out0),
     .PE_in3(PE04_out1),

     .PE_out0(PE154_out0),
     .PE_out1(PE154_out1),
     .PE_out2(PE154_out2),
     .PE_out3(PE154_out3)
       );

PE PE155(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE154_out2),
     .PE_in1(PE145_out3),
     .PE_in2(PE156_out0),
     .PE_in3(PE05_out1),

     .PE_out0(PE155_out0),
     .PE_out1(PE155_out1),
     .PE_out2(PE155_out2),
     .PE_out3(PE155_out3)
       );

PE PE156(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE155_out2),
     .PE_in1(PE146_out3),
     .PE_in2(PE157_out0),
     .PE_in3(PE06_out1),

     .PE_out0(PE156_out0),
     .PE_out1(PE156_out1),
     .PE_out2(PE156_out2),
     .PE_out3(PE156_out3)
       );

PE PE157(
     .clk(clk),
     .rst_n(rst_n),

     .PE_in0(PE156_out2),
     .PE_in1(PE147_out3),
     .PE_in2(PE150_out0),
     .PE_in3(PE07_out1),

     .PE_out0(PE157_out0),
     .PE_out1(PE157_out1),
     .PE_out2(PE157_out2),
     .PE_out3(PE157_out3)
       );



assign data_out0=PE00_out0;
assign data_out1=PE01_out0;
assign data_out2=PE02_out0;
assign data_out3=PE03_out0;

endmodule

