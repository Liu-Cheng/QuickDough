`timescale 1 ns/1 ps 

module Torus8x8 (

    Clk,
    Resetn,

    Data0_Load,
    Data0_Store,
    Data1_Load,
    Data1_Store,
    PE_Array_Busy
);

parameter DWIDTH=32;
parameter SYS_DWIDTH=32;

input                    Clk;
input                    Resetn;

input [SYS_DWIDTH-1:0]   Data0_Load;
input [SYS_DWIDTH-1:0]   Data1_Load;
output [SYS_DWIDTH-1:0]  Data0_Store;
output [SYS_DWIDTH-1:0]  Data1_Store;

input                    PE_Array_Busy;

wire [DWIDTH-1:0]        PE00_Out0;
wire [DWIDTH-1:0]        PE00_Out1;
wire [DWIDTH-1:0]        PE00_Out2;
wire [DWIDTH-1:0]        PE00_Out3;

wire [DWIDTH-1:0]        PE01_Out0;
wire [DWIDTH-1:0]        PE01_Out1;
wire [DWIDTH-1:0]        PE01_Out2;
wire [DWIDTH-1:0]        PE01_Out3;

wire [DWIDTH-1:0]        PE02_Out0;
wire [DWIDTH-1:0]        PE02_Out1;
wire [DWIDTH-1:0]        PE02_Out2;
wire [DWIDTH-1:0]        PE02_Out3;

wire [DWIDTH-1:0]        PE03_Out0;
wire [DWIDTH-1:0]        PE03_Out1;
wire [DWIDTH-1:0]        PE03_Out2;
wire [DWIDTH-1:0]        PE03_Out3;

wire [DWIDTH-1:0]        PE04_Out0;
wire [DWIDTH-1:0]        PE04_Out1;
wire [DWIDTH-1:0]        PE04_Out2;
wire [DWIDTH-1:0]        PE04_Out3;

wire [DWIDTH-1:0]        PE05_Out0;
wire [DWIDTH-1:0]        PE05_Out1;
wire [DWIDTH-1:0]        PE05_Out2;
wire [DWIDTH-1:0]        PE05_Out3;

wire [DWIDTH-1:0]        PE06_Out0;
wire [DWIDTH-1:0]        PE06_Out1;
wire [DWIDTH-1:0]        PE06_Out2;
wire [DWIDTH-1:0]        PE06_Out3;

wire [DWIDTH-1:0]        PE07_Out0;
wire [DWIDTH-1:0]        PE07_Out1;
wire [DWIDTH-1:0]        PE07_Out2;
wire [DWIDTH-1:0]        PE07_Out3;

wire [DWIDTH-1:0]        PE10_Out0;
wire [DWIDTH-1:0]        PE10_Out1;
wire [DWIDTH-1:0]        PE10_Out2;
wire [DWIDTH-1:0]        PE10_Out3;

wire [DWIDTH-1:0]        PE11_Out0;
wire [DWIDTH-1:0]        PE11_Out1;
wire [DWIDTH-1:0]        PE11_Out2;
wire [DWIDTH-1:0]        PE11_Out3;

wire [DWIDTH-1:0]        PE12_Out0;
wire [DWIDTH-1:0]        PE12_Out1;
wire [DWIDTH-1:0]        PE12_Out2;
wire [DWIDTH-1:0]        PE12_Out3;

wire [DWIDTH-1:0]        PE13_Out0;
wire [DWIDTH-1:0]        PE13_Out1;
wire [DWIDTH-1:0]        PE13_Out2;
wire [DWIDTH-1:0]        PE13_Out3;

wire [DWIDTH-1:0]        PE14_Out0;
wire [DWIDTH-1:0]        PE14_Out1;
wire [DWIDTH-1:0]        PE14_Out2;
wire [DWIDTH-1:0]        PE14_Out3;

wire [DWIDTH-1:0]        PE15_Out0;
wire [DWIDTH-1:0]        PE15_Out1;
wire [DWIDTH-1:0]        PE15_Out2;
wire [DWIDTH-1:0]        PE15_Out3;

wire [DWIDTH-1:0]        PE16_Out0;
wire [DWIDTH-1:0]        PE16_Out1;
wire [DWIDTH-1:0]        PE16_Out2;
wire [DWIDTH-1:0]        PE16_Out3;

wire [DWIDTH-1:0]        PE17_Out0;
wire [DWIDTH-1:0]        PE17_Out1;
wire [DWIDTH-1:0]        PE17_Out2;
wire [DWIDTH-1:0]        PE17_Out3;

wire [DWIDTH-1:0]        PE20_Out0;
wire [DWIDTH-1:0]        PE20_Out1;
wire [DWIDTH-1:0]        PE20_Out2;
wire [DWIDTH-1:0]        PE20_Out3;

wire [DWIDTH-1:0]        PE21_Out0;
wire [DWIDTH-1:0]        PE21_Out1;
wire [DWIDTH-1:0]        PE21_Out2;
wire [DWIDTH-1:0]        PE21_Out3;

wire [DWIDTH-1:0]        PE22_Out0;
wire [DWIDTH-1:0]        PE22_Out1;
wire [DWIDTH-1:0]        PE22_Out2;
wire [DWIDTH-1:0]        PE22_Out3;

wire [DWIDTH-1:0]        PE23_Out0;
wire [DWIDTH-1:0]        PE23_Out1;
wire [DWIDTH-1:0]        PE23_Out2;
wire [DWIDTH-1:0]        PE23_Out3;

wire [DWIDTH-1:0]        PE24_Out0;
wire [DWIDTH-1:0]        PE24_Out1;
wire [DWIDTH-1:0]        PE24_Out2;
wire [DWIDTH-1:0]        PE24_Out3;

wire [DWIDTH-1:0]        PE25_Out0;
wire [DWIDTH-1:0]        PE25_Out1;
wire [DWIDTH-1:0]        PE25_Out2;
wire [DWIDTH-1:0]        PE25_Out3;

wire [DWIDTH-1:0]        PE26_Out0;
wire [DWIDTH-1:0]        PE26_Out1;
wire [DWIDTH-1:0]        PE26_Out2;
wire [DWIDTH-1:0]        PE26_Out3;

wire [DWIDTH-1:0]        PE27_Out0;
wire [DWIDTH-1:0]        PE27_Out1;
wire [DWIDTH-1:0]        PE27_Out2;
wire [DWIDTH-1:0]        PE27_Out3;

wire [DWIDTH-1:0]        PE30_Out0;
wire [DWIDTH-1:0]        PE30_Out1;
wire [DWIDTH-1:0]        PE30_Out2;
wire [DWIDTH-1:0]        PE30_Out3;

wire [DWIDTH-1:0]        PE31_Out0;
wire [DWIDTH-1:0]        PE31_Out1;
wire [DWIDTH-1:0]        PE31_Out2;
wire [DWIDTH-1:0]        PE31_Out3;

wire [DWIDTH-1:0]        PE32_Out0;
wire [DWIDTH-1:0]        PE32_Out1;
wire [DWIDTH-1:0]        PE32_Out2;
wire [DWIDTH-1:0]        PE32_Out3;

wire [DWIDTH-1:0]        PE33_Out0;
wire [DWIDTH-1:0]        PE33_Out1;
wire [DWIDTH-1:0]        PE33_Out2;
wire [DWIDTH-1:0]        PE33_Out3;

wire [DWIDTH-1:0]        PE34_Out0;
wire [DWIDTH-1:0]        PE34_Out1;
wire [DWIDTH-1:0]        PE34_Out2;
wire [DWIDTH-1:0]        PE34_Out3;

wire [DWIDTH-1:0]        PE35_Out0;
wire [DWIDTH-1:0]        PE35_Out1;
wire [DWIDTH-1:0]        PE35_Out2;
wire [DWIDTH-1:0]        PE35_Out3;

wire [DWIDTH-1:0]        PE36_Out0;
wire [DWIDTH-1:0]        PE36_Out1;
wire [DWIDTH-1:0]        PE36_Out2;
wire [DWIDTH-1:0]        PE36_Out3;

wire [DWIDTH-1:0]        PE37_Out0;
wire [DWIDTH-1:0]        PE37_Out1;
wire [DWIDTH-1:0]        PE37_Out2;
wire [DWIDTH-1:0]        PE37_Out3;

wire [DWIDTH-1:0]        PE40_Out0;
wire [DWIDTH-1:0]        PE40_Out1;
wire [DWIDTH-1:0]        PE40_Out2;
wire [DWIDTH-1:0]        PE40_Out3;

wire [DWIDTH-1:0]        PE41_Out0;
wire [DWIDTH-1:0]        PE41_Out1;
wire [DWIDTH-1:0]        PE41_Out2;
wire [DWIDTH-1:0]        PE41_Out3;

wire [DWIDTH-1:0]        PE42_Out0;
wire [DWIDTH-1:0]        PE42_Out1;
wire [DWIDTH-1:0]        PE42_Out2;
wire [DWIDTH-1:0]        PE42_Out3;

wire [DWIDTH-1:0]        PE43_Out0;
wire [DWIDTH-1:0]        PE43_Out1;
wire [DWIDTH-1:0]        PE43_Out2;
wire [DWIDTH-1:0]        PE43_Out3;

wire [DWIDTH-1:0]        PE44_Out0;
wire [DWIDTH-1:0]        PE44_Out1;
wire [DWIDTH-1:0]        PE44_Out2;
wire [DWIDTH-1:0]        PE44_Out3;

wire [DWIDTH-1:0]        PE45_Out0;
wire [DWIDTH-1:0]        PE45_Out1;
wire [DWIDTH-1:0]        PE45_Out2;
wire [DWIDTH-1:0]        PE45_Out3;

wire [DWIDTH-1:0]        PE46_Out0;
wire [DWIDTH-1:0]        PE46_Out1;
wire [DWIDTH-1:0]        PE46_Out2;
wire [DWIDTH-1:0]        PE46_Out3;

wire [DWIDTH-1:0]        PE47_Out0;
wire [DWIDTH-1:0]        PE47_Out1;
wire [DWIDTH-1:0]        PE47_Out2;
wire [DWIDTH-1:0]        PE47_Out3;

wire [DWIDTH-1:0]        PE50_Out0;
wire [DWIDTH-1:0]        PE50_Out1;
wire [DWIDTH-1:0]        PE50_Out2;
wire [DWIDTH-1:0]        PE50_Out3;

wire [DWIDTH-1:0]        PE51_Out0;
wire [DWIDTH-1:0]        PE51_Out1;
wire [DWIDTH-1:0]        PE51_Out2;
wire [DWIDTH-1:0]        PE51_Out3;

wire [DWIDTH-1:0]        PE52_Out0;
wire [DWIDTH-1:0]        PE52_Out1;
wire [DWIDTH-1:0]        PE52_Out2;
wire [DWIDTH-1:0]        PE52_Out3;

wire [DWIDTH-1:0]        PE53_Out0;
wire [DWIDTH-1:0]        PE53_Out1;
wire [DWIDTH-1:0]        PE53_Out2;
wire [DWIDTH-1:0]        PE53_Out3;

wire [DWIDTH-1:0]        PE54_Out0;
wire [DWIDTH-1:0]        PE54_Out1;
wire [DWIDTH-1:0]        PE54_Out2;
wire [DWIDTH-1:0]        PE54_Out3;

wire [DWIDTH-1:0]        PE55_Out0;
wire [DWIDTH-1:0]        PE55_Out1;
wire [DWIDTH-1:0]        PE55_Out2;
wire [DWIDTH-1:0]        PE55_Out3;

wire [DWIDTH-1:0]        PE56_Out0;
wire [DWIDTH-1:0]        PE56_Out1;
wire [DWIDTH-1:0]        PE56_Out2;
wire [DWIDTH-1:0]        PE56_Out3;

wire [DWIDTH-1:0]        PE57_Out0;
wire [DWIDTH-1:0]        PE57_Out1;
wire [DWIDTH-1:0]        PE57_Out2;
wire [DWIDTH-1:0]        PE57_Out3;

wire [DWIDTH-1:0]        PE60_Out0;
wire [DWIDTH-1:0]        PE60_Out1;
wire [DWIDTH-1:0]        PE60_Out2;
wire [DWIDTH-1:0]        PE60_Out3;

wire [DWIDTH-1:0]        PE61_Out0;
wire [DWIDTH-1:0]        PE61_Out1;
wire [DWIDTH-1:0]        PE61_Out2;
wire [DWIDTH-1:0]        PE61_Out3;

wire [DWIDTH-1:0]        PE62_Out0;
wire [DWIDTH-1:0]        PE62_Out1;
wire [DWIDTH-1:0]        PE62_Out2;
wire [DWIDTH-1:0]        PE62_Out3;

wire [DWIDTH-1:0]        PE63_Out0;
wire [DWIDTH-1:0]        PE63_Out1;
wire [DWIDTH-1:0]        PE63_Out2;
wire [DWIDTH-1:0]        PE63_Out3;

wire [DWIDTH-1:0]        PE64_Out0;
wire [DWIDTH-1:0]        PE64_Out1;
wire [DWIDTH-1:0]        PE64_Out2;
wire [DWIDTH-1:0]        PE64_Out3;

wire [DWIDTH-1:0]        PE65_Out0;
wire [DWIDTH-1:0]        PE65_Out1;
wire [DWIDTH-1:0]        PE65_Out2;
wire [DWIDTH-1:0]        PE65_Out3;

wire [DWIDTH-1:0]        PE66_Out0;
wire [DWIDTH-1:0]        PE66_Out1;
wire [DWIDTH-1:0]        PE66_Out2;
wire [DWIDTH-1:0]        PE66_Out3;

wire [DWIDTH-1:0]        PE67_Out0;
wire [DWIDTH-1:0]        PE67_Out1;
wire [DWIDTH-1:0]        PE67_Out2;
wire [DWIDTH-1:0]        PE67_Out3;

wire [DWIDTH-1:0]        PE70_Out0;
wire [DWIDTH-1:0]        PE70_Out1;
wire [DWIDTH-1:0]        PE70_Out2;
wire [DWIDTH-1:0]        PE70_Out3;

wire [DWIDTH-1:0]        PE71_Out0;
wire [DWIDTH-1:0]        PE71_Out1;
wire [DWIDTH-1:0]        PE71_Out2;
wire [DWIDTH-1:0]        PE71_Out3;

wire [DWIDTH-1:0]        PE72_Out0;
wire [DWIDTH-1:0]        PE72_Out1;
wire [DWIDTH-1:0]        PE72_Out2;
wire [DWIDTH-1:0]        PE72_Out3;

wire [DWIDTH-1:0]        PE73_Out0;
wire [DWIDTH-1:0]        PE73_Out1;
wire [DWIDTH-1:0]        PE73_Out2;
wire [DWIDTH-1:0]        PE73_Out3;

wire [DWIDTH-1:0]        PE74_Out0;
wire [DWIDTH-1:0]        PE74_Out1;
wire [DWIDTH-1:0]        PE74_Out2;
wire [DWIDTH-1:0]        PE74_Out3;

wire [DWIDTH-1:0]        PE75_Out0;
wire [DWIDTH-1:0]        PE75_Out1;
wire [DWIDTH-1:0]        PE75_Out2;
wire [DWIDTH-1:0]        PE75_Out3;

wire [DWIDTH-1:0]        PE76_Out0;
wire [DWIDTH-1:0]        PE76_Out1;
wire [DWIDTH-1:0]        PE76_Out2;
wire [DWIDTH-1:0]        PE76_Out3;

wire [DWIDTH-1:0]        PE77_Out0;
wire [DWIDTH-1:0]        PE77_Out1;
wire [DWIDTH-1:0]        PE77_Out2;
wire [DWIDTH-1:0]        PE77_Out3;

PEIO PE00(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE07_Out2),
    .PE_In1(PE70_Out3),
    .PE_In2(PE01_Out0),
    .PE_In3(PE10_Out1),
    .PE_Out0(PE00_Out0),
    .PE_Out1(PE00_Out1),
    .PE_Out2(PE00_Out2),
    .PE_Out3(PE00_Out3),

    .PE_Load(Data0_Load),
    .PE_Store(Data0_Store),
    .PE_Array_Busy(PE_Array_Busy)

);
PEIO PE01(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE00_Out2),
    .PE_In1(PE71_Out3),
    .PE_In2(PE02_Out0),
    .PE_In3(PE11_Out1),
    .PE_Out0(PE01_Out0),
    .PE_Out1(PE01_Out1),
    .PE_Out2(PE01_Out2),
    .PE_Out3(PE01_Out3),

    .PE_Load(Data1_Load),
    .PE_Store(Data1_Store),
    .PE_Array_Busy(PE_Array_Busy)

);
PE PE02(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE01_Out2),
    .PE_In1(PE72_Out3),
    .PE_In2(PE03_Out0),
    .PE_In3(PE12_Out1),
    .PE_Out0(PE02_Out0),
    .PE_Out1(PE02_Out1),
    .PE_Out2(PE02_Out2),
    .PE_Out3(PE02_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE03(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE02_Out2),
    .PE_In1(PE73_Out3),
    .PE_In2(PE04_Out0),
    .PE_In3(PE13_Out1),
    .PE_Out0(PE03_Out0),
    .PE_Out1(PE03_Out1),
    .PE_Out2(PE03_Out2),
    .PE_Out3(PE03_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE04(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE03_Out2),
    .PE_In1(PE74_Out3),
    .PE_In2(PE05_Out0),
    .PE_In3(PE14_Out1),
    .PE_Out0(PE04_Out0),
    .PE_Out1(PE04_Out1),
    .PE_Out2(PE04_Out2),
    .PE_Out3(PE04_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE05(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE04_Out2),
    .PE_In1(PE75_Out3),
    .PE_In2(PE06_Out0),
    .PE_In3(PE15_Out1),
    .PE_Out0(PE05_Out0),
    .PE_Out1(PE05_Out1),
    .PE_Out2(PE05_Out2),
    .PE_Out3(PE05_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE06(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE05_Out2),
    .PE_In1(PE76_Out3),
    .PE_In2(PE07_Out0),
    .PE_In3(PE16_Out1),
    .PE_Out0(PE06_Out0),
    .PE_Out1(PE06_Out1),
    .PE_Out2(PE06_Out2),
    .PE_Out3(PE06_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE07(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE06_Out2),
    .PE_In1(PE77_Out3),
    .PE_In2(PE00_Out0),
    .PE_In3(PE17_Out1),
    .PE_Out0(PE07_Out0),
    .PE_Out1(PE07_Out1),
    .PE_Out2(PE07_Out2),
    .PE_Out3(PE07_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE10(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE17_Out2),
    .PE_In1(PE00_Out3),
    .PE_In2(PE11_Out0),
    .PE_In3(PE20_Out1),
    .PE_Out0(PE10_Out0),
    .PE_Out1(PE10_Out1),
    .PE_Out2(PE10_Out2),
    .PE_Out3(PE10_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE11(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE10_Out2),
    .PE_In1(PE01_Out3),
    .PE_In2(PE12_Out0),
    .PE_In3(PE21_Out1),
    .PE_Out0(PE11_Out0),
    .PE_Out1(PE11_Out1),
    .PE_Out2(PE11_Out2),
    .PE_Out3(PE11_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE12(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE11_Out2),
    .PE_In1(PE02_Out3),
    .PE_In2(PE13_Out0),
    .PE_In3(PE22_Out1),
    .PE_Out0(PE12_Out0),
    .PE_Out1(PE12_Out1),
    .PE_Out2(PE12_Out2),
    .PE_Out3(PE12_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE13(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE12_Out2),
    .PE_In1(PE03_Out3),
    .PE_In2(PE14_Out0),
    .PE_In3(PE23_Out1),
    .PE_Out0(PE13_Out0),
    .PE_Out1(PE13_Out1),
    .PE_Out2(PE13_Out2),
    .PE_Out3(PE13_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE14(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE13_Out2),
    .PE_In1(PE04_Out3),
    .PE_In2(PE15_Out0),
    .PE_In3(PE24_Out1),
    .PE_Out0(PE14_Out0),
    .PE_Out1(PE14_Out1),
    .PE_Out2(PE14_Out2),
    .PE_Out3(PE14_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE15(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE14_Out2),
    .PE_In1(PE05_Out3),
    .PE_In2(PE16_Out0),
    .PE_In3(PE25_Out1),
    .PE_Out0(PE15_Out0),
    .PE_Out1(PE15_Out1),
    .PE_Out2(PE15_Out2),
    .PE_Out3(PE15_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE16(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE15_Out2),
    .PE_In1(PE06_Out3),
    .PE_In2(PE17_Out0),
    .PE_In3(PE26_Out1),
    .PE_Out0(PE16_Out0),
    .PE_Out1(PE16_Out1),
    .PE_Out2(PE16_Out2),
    .PE_Out3(PE16_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE17(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE16_Out2),
    .PE_In1(PE07_Out3),
    .PE_In2(PE10_Out0),
    .PE_In3(PE27_Out1),
    .PE_Out0(PE17_Out0),
    .PE_Out1(PE17_Out1),
    .PE_Out2(PE17_Out2),
    .PE_Out3(PE17_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE20(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE27_Out2),
    .PE_In1(PE10_Out3),
    .PE_In2(PE21_Out0),
    .PE_In3(PE30_Out1),
    .PE_Out0(PE20_Out0),
    .PE_Out1(PE20_Out1),
    .PE_Out2(PE20_Out2),
    .PE_Out3(PE20_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE21(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE20_Out2),
    .PE_In1(PE11_Out3),
    .PE_In2(PE22_Out0),
    .PE_In3(PE31_Out1),
    .PE_Out0(PE21_Out0),
    .PE_Out1(PE21_Out1),
    .PE_Out2(PE21_Out2),
    .PE_Out3(PE21_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE22(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE21_Out2),
    .PE_In1(PE12_Out3),
    .PE_In2(PE23_Out0),
    .PE_In3(PE32_Out1),
    .PE_Out0(PE22_Out0),
    .PE_Out1(PE22_Out1),
    .PE_Out2(PE22_Out2),
    .PE_Out3(PE22_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE23(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE22_Out2),
    .PE_In1(PE13_Out3),
    .PE_In2(PE24_Out0),
    .PE_In3(PE33_Out1),
    .PE_Out0(PE23_Out0),
    .PE_Out1(PE23_Out1),
    .PE_Out2(PE23_Out2),
    .PE_Out3(PE23_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE24(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE23_Out2),
    .PE_In1(PE14_Out3),
    .PE_In2(PE25_Out0),
    .PE_In3(PE34_Out1),
    .PE_Out0(PE24_Out0),
    .PE_Out1(PE24_Out1),
    .PE_Out2(PE24_Out2),
    .PE_Out3(PE24_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE25(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE24_Out2),
    .PE_In1(PE15_Out3),
    .PE_In2(PE26_Out0),
    .PE_In3(PE35_Out1),
    .PE_Out0(PE25_Out0),
    .PE_Out1(PE25_Out1),
    .PE_Out2(PE25_Out2),
    .PE_Out3(PE25_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE26(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE25_Out2),
    .PE_In1(PE16_Out3),
    .PE_In2(PE27_Out0),
    .PE_In3(PE36_Out1),
    .PE_Out0(PE26_Out0),
    .PE_Out1(PE26_Out1),
    .PE_Out2(PE26_Out2),
    .PE_Out3(PE26_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE27(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE26_Out2),
    .PE_In1(PE17_Out3),
    .PE_In2(PE20_Out0),
    .PE_In3(PE37_Out1),
    .PE_Out0(PE27_Out0),
    .PE_Out1(PE27_Out1),
    .PE_Out2(PE27_Out2),
    .PE_Out3(PE27_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE30(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE37_Out2),
    .PE_In1(PE20_Out3),
    .PE_In2(PE31_Out0),
    .PE_In3(PE40_Out1),
    .PE_Out0(PE30_Out0),
    .PE_Out1(PE30_Out1),
    .PE_Out2(PE30_Out2),
    .PE_Out3(PE30_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE31(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE30_Out2),
    .PE_In1(PE21_Out3),
    .PE_In2(PE32_Out0),
    .PE_In3(PE41_Out1),
    .PE_Out0(PE31_Out0),
    .PE_Out1(PE31_Out1),
    .PE_Out2(PE31_Out2),
    .PE_Out3(PE31_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE32(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE31_Out2),
    .PE_In1(PE22_Out3),
    .PE_In2(PE33_Out0),
    .PE_In3(PE42_Out1),
    .PE_Out0(PE32_Out0),
    .PE_Out1(PE32_Out1),
    .PE_Out2(PE32_Out2),
    .PE_Out3(PE32_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE33(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE32_Out2),
    .PE_In1(PE23_Out3),
    .PE_In2(PE34_Out0),
    .PE_In3(PE43_Out1),
    .PE_Out0(PE33_Out0),
    .PE_Out1(PE33_Out1),
    .PE_Out2(PE33_Out2),
    .PE_Out3(PE33_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE34(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE33_Out2),
    .PE_In1(PE24_Out3),
    .PE_In2(PE35_Out0),
    .PE_In3(PE44_Out1),
    .PE_Out0(PE34_Out0),
    .PE_Out1(PE34_Out1),
    .PE_Out2(PE34_Out2),
    .PE_Out3(PE34_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE35(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE34_Out2),
    .PE_In1(PE25_Out3),
    .PE_In2(PE36_Out0),
    .PE_In3(PE45_Out1),
    .PE_Out0(PE35_Out0),
    .PE_Out1(PE35_Out1),
    .PE_Out2(PE35_Out2),
    .PE_Out3(PE35_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE36(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE35_Out2),
    .PE_In1(PE26_Out3),
    .PE_In2(PE37_Out0),
    .PE_In3(PE46_Out1),
    .PE_Out0(PE36_Out0),
    .PE_Out1(PE36_Out1),
    .PE_Out2(PE36_Out2),
    .PE_Out3(PE36_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE37(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE36_Out2),
    .PE_In1(PE27_Out3),
    .PE_In2(PE30_Out0),
    .PE_In3(PE47_Out1),
    .PE_Out0(PE37_Out0),
    .PE_Out1(PE37_Out1),
    .PE_Out2(PE37_Out2),
    .PE_Out3(PE37_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE40(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE47_Out2),
    .PE_In1(PE30_Out3),
    .PE_In2(PE41_Out0),
    .PE_In3(PE50_Out1),
    .PE_Out0(PE40_Out0),
    .PE_Out1(PE40_Out1),
    .PE_Out2(PE40_Out2),
    .PE_Out3(PE40_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE41(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE40_Out2),
    .PE_In1(PE31_Out3),
    .PE_In2(PE42_Out0),
    .PE_In3(PE51_Out1),
    .PE_Out0(PE41_Out0),
    .PE_Out1(PE41_Out1),
    .PE_Out2(PE41_Out2),
    .PE_Out3(PE41_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE42(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE41_Out2),
    .PE_In1(PE32_Out3),
    .PE_In2(PE43_Out0),
    .PE_In3(PE52_Out1),
    .PE_Out0(PE42_Out0),
    .PE_Out1(PE42_Out1),
    .PE_Out2(PE42_Out2),
    .PE_Out3(PE42_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE43(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE42_Out2),
    .PE_In1(PE33_Out3),
    .PE_In2(PE44_Out0),
    .PE_In3(PE53_Out1),
    .PE_Out0(PE43_Out0),
    .PE_Out1(PE43_Out1),
    .PE_Out2(PE43_Out2),
    .PE_Out3(PE43_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE44(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE43_Out2),
    .PE_In1(PE34_Out3),
    .PE_In2(PE45_Out0),
    .PE_In3(PE54_Out1),
    .PE_Out0(PE44_Out0),
    .PE_Out1(PE44_Out1),
    .PE_Out2(PE44_Out2),
    .PE_Out3(PE44_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE45(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE44_Out2),
    .PE_In1(PE35_Out3),
    .PE_In2(PE46_Out0),
    .PE_In3(PE55_Out1),
    .PE_Out0(PE45_Out0),
    .PE_Out1(PE45_Out1),
    .PE_Out2(PE45_Out2),
    .PE_Out3(PE45_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE46(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE45_Out2),
    .PE_In1(PE36_Out3),
    .PE_In2(PE47_Out0),
    .PE_In3(PE56_Out1),
    .PE_Out0(PE46_Out0),
    .PE_Out1(PE46_Out1),
    .PE_Out2(PE46_Out2),
    .PE_Out3(PE46_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE47(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE46_Out2),
    .PE_In1(PE37_Out3),
    .PE_In2(PE40_Out0),
    .PE_In3(PE57_Out1),
    .PE_Out0(PE47_Out0),
    .PE_Out1(PE47_Out1),
    .PE_Out2(PE47_Out2),
    .PE_Out3(PE47_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE50(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE57_Out2),
    .PE_In1(PE40_Out3),
    .PE_In2(PE51_Out0),
    .PE_In3(PE60_Out1),
    .PE_Out0(PE50_Out0),
    .PE_Out1(PE50_Out1),
    .PE_Out2(PE50_Out2),
    .PE_Out3(PE50_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE51(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE50_Out2),
    .PE_In1(PE41_Out3),
    .PE_In2(PE52_Out0),
    .PE_In3(PE61_Out1),
    .PE_Out0(PE51_Out0),
    .PE_Out1(PE51_Out1),
    .PE_Out2(PE51_Out2),
    .PE_Out3(PE51_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE52(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE51_Out2),
    .PE_In1(PE42_Out3),
    .PE_In2(PE53_Out0),
    .PE_In3(PE62_Out1),
    .PE_Out0(PE52_Out0),
    .PE_Out1(PE52_Out1),
    .PE_Out2(PE52_Out2),
    .PE_Out3(PE52_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE53(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE52_Out2),
    .PE_In1(PE43_Out3),
    .PE_In2(PE54_Out0),
    .PE_In3(PE63_Out1),
    .PE_Out0(PE53_Out0),
    .PE_Out1(PE53_Out1),
    .PE_Out2(PE53_Out2),
    .PE_Out3(PE53_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE54(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE53_Out2),
    .PE_In1(PE44_Out3),
    .PE_In2(PE55_Out0),
    .PE_In3(PE64_Out1),
    .PE_Out0(PE54_Out0),
    .PE_Out1(PE54_Out1),
    .PE_Out2(PE54_Out2),
    .PE_Out3(PE54_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE55(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE54_Out2),
    .PE_In1(PE45_Out3),
    .PE_In2(PE56_Out0),
    .PE_In3(PE65_Out1),
    .PE_Out0(PE55_Out0),
    .PE_Out1(PE55_Out1),
    .PE_Out2(PE55_Out2),
    .PE_Out3(PE55_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE56(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE55_Out2),
    .PE_In1(PE46_Out3),
    .PE_In2(PE57_Out0),
    .PE_In3(PE66_Out1),
    .PE_Out0(PE56_Out0),
    .PE_Out1(PE56_Out1),
    .PE_Out2(PE56_Out2),
    .PE_Out3(PE56_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE57(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE56_Out2),
    .PE_In1(PE47_Out3),
    .PE_In2(PE50_Out0),
    .PE_In3(PE67_Out1),
    .PE_Out0(PE57_Out0),
    .PE_Out1(PE57_Out1),
    .PE_Out2(PE57_Out2),
    .PE_Out3(PE57_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE60(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE67_Out2),
    .PE_In1(PE50_Out3),
    .PE_In2(PE61_Out0),
    .PE_In3(PE70_Out1),
    .PE_Out0(PE60_Out0),
    .PE_Out1(PE60_Out1),
    .PE_Out2(PE60_Out2),
    .PE_Out3(PE60_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE61(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE60_Out2),
    .PE_In1(PE51_Out3),
    .PE_In2(PE62_Out0),
    .PE_In3(PE71_Out1),
    .PE_Out0(PE61_Out0),
    .PE_Out1(PE61_Out1),
    .PE_Out2(PE61_Out2),
    .PE_Out3(PE61_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE62(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE61_Out2),
    .PE_In1(PE52_Out3),
    .PE_In2(PE63_Out0),
    .PE_In3(PE72_Out1),
    .PE_Out0(PE62_Out0),
    .PE_Out1(PE62_Out1),
    .PE_Out2(PE62_Out2),
    .PE_Out3(PE62_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE63(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE62_Out2),
    .PE_In1(PE53_Out3),
    .PE_In2(PE64_Out0),
    .PE_In3(PE73_Out1),
    .PE_Out0(PE63_Out0),
    .PE_Out1(PE63_Out1),
    .PE_Out2(PE63_Out2),
    .PE_Out3(PE63_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE64(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE63_Out2),
    .PE_In1(PE54_Out3),
    .PE_In2(PE65_Out0),
    .PE_In3(PE74_Out1),
    .PE_Out0(PE64_Out0),
    .PE_Out1(PE64_Out1),
    .PE_Out2(PE64_Out2),
    .PE_Out3(PE64_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE65(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE64_Out2),
    .PE_In1(PE55_Out3),
    .PE_In2(PE66_Out0),
    .PE_In3(PE75_Out1),
    .PE_Out0(PE65_Out0),
    .PE_Out1(PE65_Out1),
    .PE_Out2(PE65_Out2),
    .PE_Out3(PE65_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE66(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE65_Out2),
    .PE_In1(PE56_Out3),
    .PE_In2(PE67_Out0),
    .PE_In3(PE76_Out1),
    .PE_Out0(PE66_Out0),
    .PE_Out1(PE66_Out1),
    .PE_Out2(PE66_Out2),
    .PE_Out3(PE66_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE67(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE66_Out2),
    .PE_In1(PE57_Out3),
    .PE_In2(PE60_Out0),
    .PE_In3(PE77_Out1),
    .PE_Out0(PE67_Out0),
    .PE_Out1(PE67_Out1),
    .PE_Out2(PE67_Out2),
    .PE_Out3(PE67_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE70(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE77_Out2),
    .PE_In1(PE60_Out3),
    .PE_In2(PE71_Out0),
    .PE_In3(PE00_Out1),
    .PE_Out0(PE70_Out0),
    .PE_Out1(PE70_Out1),
    .PE_Out2(PE70_Out2),
    .PE_Out3(PE70_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE71(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE70_Out2),
    .PE_In1(PE61_Out3),
    .PE_In2(PE72_Out0),
    .PE_In3(PE01_Out1),
    .PE_Out0(PE71_Out0),
    .PE_Out1(PE71_Out1),
    .PE_Out2(PE71_Out2),
    .PE_Out3(PE71_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE72(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE71_Out2),
    .PE_In1(PE62_Out3),
    .PE_In2(PE73_Out0),
    .PE_In3(PE02_Out1),
    .PE_Out0(PE72_Out0),
    .PE_Out1(PE72_Out1),
    .PE_Out2(PE72_Out2),
    .PE_Out3(PE72_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE73(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE72_Out2),
    .PE_In1(PE63_Out3),
    .PE_In2(PE74_Out0),
    .PE_In3(PE03_Out1),
    .PE_Out0(PE73_Out0),
    .PE_Out1(PE73_Out1),
    .PE_Out2(PE73_Out2),
    .PE_Out3(PE73_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE74(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE73_Out2),
    .PE_In1(PE64_Out3),
    .PE_In2(PE75_Out0),
    .PE_In3(PE04_Out1),
    .PE_Out0(PE74_Out0),
    .PE_Out1(PE74_Out1),
    .PE_Out2(PE74_Out2),
    .PE_Out3(PE74_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE75(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE74_Out2),
    .PE_In1(PE65_Out3),
    .PE_In2(PE76_Out0),
    .PE_In3(PE05_Out1),
    .PE_Out0(PE75_Out0),
    .PE_Out1(PE75_Out1),
    .PE_Out2(PE75_Out2),
    .PE_Out3(PE75_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE76(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE75_Out2),
    .PE_In1(PE66_Out3),
    .PE_In2(PE77_Out0),
    .PE_In3(PE06_Out1),
    .PE_Out0(PE76_Out0),
    .PE_Out1(PE76_Out1),
    .PE_Out2(PE76_Out2),
    .PE_Out3(PE76_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
PE PE77(
    .Clk(Clk),
    .Resetn(Resetn),

    .PE_In0(PE76_Out2),
    .PE_In1(PE67_Out3),
    .PE_In2(PE70_Out0),
    .PE_In3(PE07_Out1),
    .PE_Out0(PE77_Out0),
    .PE_Out1(PE77_Out1),
    .PE_Out2(PE77_Out2),
    .PE_Out3(PE77_Out3),

    .PE_Array_Busy(PE_Array_Busy)

);
endmodule
